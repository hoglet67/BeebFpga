`timescale 1ns / 1ns

`define p1edge posedge
`define p2edge posedge

module hp_flag_m

`include "gen_flag_v3.v"

--
--Written by GowinSynthesis
--Tool Version "V1.9.11"
--Tue Jan 28 15:02:31 2025

--Source file index table:
--file0 "\/disk1/home/dmb/atom/BeebFpga/src/gowin/tang20k/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_define.v"
--file1 "\/disk1/home/dmb/atom/BeebFpga/src/gowin/tang20k/src/fifo_sc_hs/temp/FIFO_SC/fifo_sc_hs_parameter.v"
--file2 "\/disk1/home/dmb/gowin/v1.9.11/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs.v"
--file3 "\/disk1/home/dmb/gowin/v1.9.11/IDE/ipcore/FIFO_SC_HS/data/fifo_sc_hs_top.v"
`protect begin_protected
`protect version="2.3"
`protect author="default"
`protect author_info="default"
`protect encrypt_agent="GOWIN"
`protect encrypt_agent_info="GOWIN Encrypt Version 2.3"

`protect encoding=(enctype="base64", line_length=76, bytes=256)
`protect key_keyowner="GOWIN",key_keyname="GWK2023-09",key_method="rsa"
`protect key_block
hGXaPSYxlhxkdo1xFLsABTQdEw39Y7ApKtK/OaOXEDrTpSt6v8nB5LQiJoyhoZOuNff2+ZAmsr8d
WQfl6RF0dBNsDk8gM7lQ0euXxDoxwv5wLB/u/z0VoPW8ink0fF7/XbxyllpbteAzhiEs+isQMTGq
/QX+EwPYG4JNThlOwDek1wrPHCtUK4xgOOIcECe4S/JX8F6M5e/wtJmewH7vt+odRABasSKwWgP+
nlcPKoA/NaYkN/nVeaS4LJTzzs7eg7cLiUZamV3MknMuKOACnS3T/MccYZRr9hytlYLh7iHX8M56
fHy5ir7H0n5UJOe9kA1ZYg4HaSou7FCYPAr4FA==

`protect encoding=(enctype="base64", line_length=76, bytes=15760)
`protect data_keyowner="default-ip-vendor"
`protect data_keyname="default-ip-key"
`protect data_method="aes128-cfb"
`protect data_block
wKANodWVVo/5LT/bAOBJqeTurWaC0J0tUryTvDvvHTfKoaedmEy/r4OBq7TcNhC0Nt1HmGZ1opqc
0+H0r5K8LNX4C8fpYcX30fR5AigsqbL8sizyPYbXMO9wzfdiO8SYrjwFqAdVBvu5ynFbv8z8rqre
ZKbsYcRTrbDXCJHEHyXrmlf6wlFw+m6EOswoPLC9EEN5/HNNENSQOf81XT+MTsmUiXx+MfIC8Gts
Bs7JJc+8pcihZstnWAiFk/AkYLLqH6qVX+4IXxjy2OT7PbKZQxcFsTuGyr3GydLF8DVvXqw295xQ
cq1VMsAesJt5rS6BLu3OzlC/qRt3yVxbC19xonNHcgpN8M3KjnmfeIhL3LP5LRn86FHj9RuWo0vs
pW+wz5ZyrUqU3XUXIg//0uAGuGMprK+EuFVBflbuf1zZpL/+1cCPoD8yCZkJpIC7m60+iODoI3nA
YG/JrVMTBrA9Aq0kMk9Tf7weIj2Npcsk+Qgue3z/xWSa9S8bWGbB53V/1d//kq6kvQSDZirYGjrY
9/6G6Av0B/al3fnUT5tSMRXz8cAAjbTozTJ7d1YtXGn+vHTZl74LaPHxpPtjslSxwJBfWxb6bVFZ
o2UtLz+rTK6cR4N/9k9Ykf3BPxaV5bHV6zwtQSqlAhYy1ArRSsGQ2ktQdgBDZnh4JiEzbMCtqZo6
0ihrJWKFGARoya5TXIqvDsIQQUXYh94864wqhUie8QlVCVSHHZKv/IURAl41ggcQs/HXeT1shKZZ
bfuqus27v+JmZ2iAtzfVtI89Q53O1guoyRmo3ce02gvmLo7EkpyLBgKPD2TwC3mPsa2eDTDXlu7r
j/hHpTQwwxlRrMTkqXCyuZCEgb6pUAbuDi8jox2PIp3Wv4Rb1o3t3xQ9h+/na09L5UppyAnaWAt7
k0Fi+4SbKJbD0jzqiO6mfYfAEQhXgn7QIr/3IIUwwH05TUTeaP+p7Rdcvm6R6HnCq8x5Wf3Rw/YX
xS2wyw4rqwUQuCQvOMZk3S56nPFET2V607bGW2l5PoPHKP+QmJQGuYOaZpEZq0//pGOl+W4shmvb
nV7BGA1zckiMj2/m5lXovR/XSVa+kBtmWoRW/BzctDLKOBPjGzY9grepLajBeHnNMfNsW6JY9ofc
YWFpzD5mhYYPX7O5AKhafmNS2O2nFvM1Lb+JtM8dn77MiKHU5maGP15ylTp/XZg0USBRbWl6U6KE
TChz9WWRZflPVbAMnKt0o2uroJ9GvMB+PHwqGjUQN+D+8P+nsreRAP82k0dnRoIjXDWImVO6g93E
I+m6eo1raY3DIG89zkwlpIC0Cbr4yzwb894xbI/tjZwGev+7ISr6rYI6yGatkni8MUtMpvwFgpov
Vbftu62te6Mk+aq+zL5RvgJBm2z+wF5MFlsYiTTuSnGd9fOEYZRJtOvN6WaqEh8qmR1TiTmBk+HJ
/7sgk07ISxkRwbYsExR1k64U25SysKz4BalPmJjLWKycFLmA7LJY12ggbuRJW5c0XQYpg/eq6YHt
x21YgeOPVczpVTQAI3oZbP1WxW4JnAmZFiEv0Z7OFfpfKtESLhmFtNDFJKkJR3stUB2ZHqiEoRAH
8wkuceGX8+fJReV4AvEc+NzNS6JB9l8GXlWv5iZkHlYMQXTchMTICPEUEx216Q+2HQzR2BddrIC3
BbAOfz6fDmO9LzYT46f7urrX86mUGN4hYQA1d9JAljOfOdx+ju0anXljW+h2aAwYoVOjhqZUJSZq
GmuR6GIYXBg8jByK2sN05Dd/ie7/WEg0hRP8K/du1kg0OoKPqDZNDAyk24iFTMO57ZAQSDXZzkOa
YwSONLXg7SAvokkkvTr8eABSZivZVD9kBoYsZ6Q2qQQphqpHA2ca8jtw1QuWSAniNJRhAquiSsc+
Br9LUPwUCcMMI+IA5rujyxf55I2aDT/BB7Ldoj6jJVB3l2+zlVGUlzW/+mZtqUr9W4dTUddD20+M
KGx1bqJyGarWdja0+K6dlh8k3YTq88afze6RiZ/0eI5pP4mTB26QkJWBjcbDHHZYccfYTC44cC8c
h8S4SzECH1dMBzCyrw3re9gXX5PgrnwwovF839/XTzam4gX3K5X8qO3BKpwGTuOSF+JBy/JLeur/
hwDnJ0bd0Noictzt43kRveVcYk75asHzjHy5O9hwedGQ54KdaUb6FIrhNiPuqC+PkrvOmuTTaGEn
D2eFwAV/3hrg4vG1oHKUtcyKWOYphRGOnFdK+ztrl17Jr8D/T0vChG2Jo69DNHpDvBDN+x+a/e7n
R564Ll2MEqkcvVAcakwOSxAUa963AmzBKijDlXI9Ka7p/XomlWwRR57Gq7LMJFx57qCadL37gQLC
8qBaMd7xge7we58VeXDXymMWu0LjuTqPNrPi1I541mhyfhqTOdI4mUwaT+20S5UkNnfYY9Ghw4vR
nNGdKcOFqWL69pET3sG1sC98OLzosedDsQeXFD7HZclZD0KVzK+aAs0uXSRp/oTPrCK69cF74WBe
bP+QC9Nkc4ujsff7I94kSPU6DO8YgMi1rMeOUOSZU3tWCvB5qSOifOiHT78LO/KiENjGfZxw6vtC
jFemGYucbqlj29drY+biGYWiSmPUd9/PLYE2DmBLTY93U9qcTsq4137AasP0iqYkfnS8FYWqSZOZ
tGkhK1iwiGF14grg5UoanXEzvsxhNv6ZqmQv23T2Ml8QVSykUdHPVZ0ViSIl4enq/6jyR9bueLVC
kDj6e3XbCiWYH3Tu5O9rK4qGu3f6FwdqP+UUknw5os5r2bem9xiXDgE736oF6bCSfQIeAq8/uvOA
e7i0LOnrTzkK7D+ZDKfpMxop29qrz8adosE4laMrNkCS5gQrZvByEYBCpSeBzpwVt5aPZIT6l//1
7Mf0n4lJqF7iU6NxFImQbrJG6QvNrp18snNxj/SC1u12lusAWZ223uBDemeGAHHwi3z7RR51O6by
42T9HMLu4Lv7FgyGHMD29e7iszvBBRar+N0aqnFYRmSeJyoncWmda6JztnuLTBLi+0zkDBxeqprC
qhfDrm+wLer5SNLiBDfd+/tzh2kih6zL/3AYQry3YkikvEnA75llu3aFi92ioJk+OyNIEX0oHn2g
0Xr/T1tVDLXlixleHwHcz3J+k/3hLxxa6eFjjsVKu+R6/633yolomjuxhOExlrmNR+xQbAItW3Nn
xO+w+J7AUhqDoYlMy9GK73A9oxWnPCPEXcS0Y6sZYmmy3B/5FGsn2xP69izutOMSdWtgi8skd2L9
0pAYHFQUz0qHy//+0OP2fwBfQ58DI+p3hekGX/br73CuHYskBE7J0LlPtrXw3KUCxFbwPaJLLR4+
PKCWm7lK/ydlGA+ce5H7v7BeQStcuCDNEdAP+U4JcYUBJBh/aZIwmbuFFG/4gKwZtgS3KYq1SlQ7
oIBVDvQ7419BGcRNApbwEmapnp607dxAsTq4XOsAfOH8uxZpjnW+nVQ0LTL40fz7HSpf4WvmP/eH
3qFSOT4PeM9LpLCZU4uRzK8+C0Ku8W22IrPhi/bIjthroF9oJFXmFXatM06cO0h3aHD5deOGY1NR
NtbXwuJEA5oF2CvMvfbTvAh1RYi+HSv+VzDB2DAhzGG5oHg6yNzy2oyo0ayi8MCQ07+iKfmnciGt
ZsXJpw/8uu/Gqvl2Gr54LuGbsDLsnLa66JuAMNdz8s7XtzMTAyeCj7lqJCi2QNZ9CdedUZPYWf6y
yC7H87lMYW0Hq+cIdJS1akReIuHQTqVeFzvBJjRQ5SeKNc9xpBuJtczETlT3Ske+/VfTGuf1X/Y4
HHLF5ludzzDSVbc6l3kmNeb/u1Qr8YUpyCw4BGY4yhgWbE+EJTJwBjBnT2JzuH+Tcyx+JQ4bff17
wmOG3e5ApXnY6ZCBIWPEmnxxNCbo95aKyiIBfmmNgsO5vs8z/jQtILTsq6+eK1iZum2wC4hcIY8I
j5P9z2UBM/qiz7LDLVcdUz6GZ2SssSfg/+ZbKfkp1WuK6LtPCI67TB+vtBW03Hl69wQvu1hYf2T+
TEzeyphWEqYHQ/iM21w07CEUs0Ovr1+gFYkYAz0DXAwmt/b6j0GTTlJZhk3olYjB84q0PhRUEJmp
fQ5T4jwUXPicDFdEWQZAJUOJ5ucR6lFK5q45JpsmYMhr80sGh5pISSBiHgmshBf+zcl/cHw+zQqm
R6dEp7RO5RE5uVOIvfV0iOWqSRXUN/hmFxdrapz9jAdNDnSWPoRIRicvLhQC7p417tHKXBUXnN9e
d0UslWvH3iaGllEJi/Fuj9RP+BkrPgSUjG0zUIeibcfUxnZXiv4oJ+0nfyGDz+vCkm83aSCNfiEp
6Ys3e2ve4P8x1N+xzTVI9Z05KhylNgW8glomu3YUybKUEvwLL9nFeI9GlMYmRdHYsb6wjbikBoog
6hmLszxhlNse0mjCtrZudVHxJeNEm0hSk6kzAV89rR8wuC/2g876JOoVYDvaLtMe9l2ohZSyrkhY
6Qi0Lss3lpukS0JaE2HSPPs6mzu6KMyba9Uzc486yFUf/KzDedVoZP1GyfslD6RrWJYIr9WQ4YKG
wYg5gzN6IVTRCbrr/ZgPlUZOrNAj+mdWOPgmXe3a7uJdUCEYOm72VhAyLfESpvPfnGmQJCPMppNs
ftIEba0PXazC92CfyvgFrDOuo/tBPvAkIs2SDS7cJhvjMayJpsLcycd566z91JZ9P2N396awQzEY
YR6fwE1LeAb6FtLIvNBxF1/4gnxv6XNbwA3M85AlhT5C2YtLwcYI/rwxXEe53+6goKF7rNqnfkrV
eC/Ks5KrG4BPzNa0Fz8XXitakZBxC0zxakAfy8eNT23sc/ShVAL+EQssV4MH5/Zo1yTNxWAgm4Ki
dW4NkvinBjRVHGC4bUMd/uZjUjpaY/L9H4AA9ZHyoTzdqrN5a7NJ6gc0UUOhE3ANi4eXjg6w0Krd
ObR7r0CN0fJFt1JCaS96XaEiH2B3IfNhnXYzZ7tWZQ6upgz+7x5Rw4nMC+VvB6Mkt3GROjZjj9xT
HT3IKOXamtvuxKO/zk2WbQnsfayqawSYzfwlDwvkIlnUte/xqByVzoD3KgPtMG+uwMK8mC34KAe1
VL5oV9Pe/PLzjPmGJkC7sD9KsSLi/ZIiPeh/4K+BYfZ1L2VKdGDXqpjF/Q7HRO0QQqbrvh3NhjNW
w2tiylN1A1+y0MgModBxz0y2LbZ81CnfgldxZF/33DjgdSYZzFNSVeFVPG2sL1iGHcfGG7q/QCGJ
IjAWtkyMMdA/lQiGXvi7qrgMCE3R9f49PoZBlHF3uaRSulCBkPpFkBVLVVN+GfCbSqiqcBizb4X7
kGZKADe9qWUVE8UViAei45aQmZZRMVxvMC77TxTKoEkWfPw+D20MSGBxsWL2xxzF1mk3uSMX+S6F
3jZR/hXyjBv5YG3N5nad6Jdw54J8ZvAXfi6KD8Ohuv60xwvuWxGATrli2rDiB0EfLeuboSbZsu09
cM7ZH47L9a9+YPe+kGgewsgMmw4KdE3o2CEXZnzpfSC4uI8UGEA9KlX7ccLFkdiq+ER0rEQqiouB
qR4uzfF7UOV9Tc9ykz+tXdaX/EPGSKMG5EEQpTaU1cU2UaKqF1Pfw4QW/QOcsKncuswjh5Bl3piD
VW5JcD2CJ8ectO6l8/FD1iE2+WHsIIUgUzUynHemGckATeqZeG/fUk/pJiuI84eHdS5pjlSnYQLf
hQsy12/Ljc2Ld4zSg5fuemXCKnhTs/YCN9u9MzniRjvoL1lG4Ve/SegIbAMqdQXXkyXXuWqVv2Kq
/1Hl9Q9WFIuhYVUcmHXPWySW8WQPQF2PPRfH9TdBNhpR6j369zLzGMODZMFIPoUEZC4b8gmBHrbf
+pC2TbyfdtS5t2mC3ErKlCiYb6pSZHTi2SO3n/f+kDbxitkIk0TUD//NcH6F5xN4VXwxCginDnHF
VK0Rbsqw9nWTcUYl6+tDT1xayHvPCrAz7dD+Aq+7tfLugyco2db0gfg6RWhJsLKNSVUQlaPgZL25
4Xct8S9bGRtfyjCYarzLjVOjlpTC1g0n6DTb/DEm6vd4lySZFHA2sfhvB6oK51gBxq6bSjtovZCR
ykLaS7pZPqan/idZeBRSgymuu5RofI0hgdhiEJiyU5F5804ChS48Q1gkczmpCu63CX+7x+It4lim
hqeUrPn87HGAza7u5/PdYE/wAQYzDkFcL+vGvs9+UaO3w7ajPaZWn4Or9CLtWp3a81SkuCwWDeXY
trosm4ZkLMpMBo4rOlslZvhFyuztfFlq2BdADJTEteZ1HaKR1zlOkGyskoC/8jgptEqLXb6fF0X/
QZYO6ogtT3G8LmucuP+7OymKacEo9zmlO3tf2mksuFrhg/56AyLWN+hjcxZQQ9CyeCZfvZxn7BDB
hEjpwxMn3SA14nDBbdYynYUHpTXOSUUcj2sq0uMd1da9rAX26qaBImX3yts/95RqyGhdLCOao6BI
9OAwiOwjHceTKXxIIWB9i+i3JzY0wcKvOWNQhTQy30+HmDCmEi4RL63tYe9eDCT2mCbvYo6CVCoR
vVQbHBmXvdBL6f4DPNsDm49TstKWd+NHnMUnxbw/fKipOZ/qCQrax8a6FwnIMFlTevjDH8GCTvU4
IEO/IJYJvZU+s+D09LKNZz/Wc8oxCfGRtdEqzA2W738LMnPSHrYzdjBmzAVn6aYql/QypGhDJV+Y
1KX8QtwjzUoGs0Y6hA6C929s616HDb+Z7Q0JoXKnFvMLkFHYmG2u2feh/Dhedckp49HvYzDZ2sFb
+A9AVgy+YzNkql3Q4Dd7zPrLIr7GNe0TjW63KHfaHWan/v2y3+Zy2DBuRt/3pNH8lOGVbmc1sqts
8d/qau25nMWTuRM+cNLPJ60drguXPDLVG9nNvmLc2kOy9FQ/A9wtT1Y6JOJcUznd7CcJgInbuB88
PkqWEnhyZWNgeB1JAiWoaaIT8dq56tfn2ofXFJGKjhUcS7aNYEUAT9Qc7JC8xTzMnJVNSF2KlvhS
NA5RMGeb8c19BzeOs8Mf6NFyJZlNTGNYIuO5ssQ/uEnuua1hoHJNh8N8XMD4Yyn/De2otdENKMLX
Y5VUsxJ0QH/lPw5JHWHmuH2L4djsMVo22JdEfO0Hs7gneuSzPWe/40dvaH9gZjB2zehiU55zM3ah
2dRuGb+LmA5gdctObbeBjANHsbCghONuWGvX/cCDzhxEt0rzIY4bgRmfjksjAlC/c5aYp7nyt4w2
zvN7gRYR9HayWAiE5kJ8a2LU6MMUcIDHWQsp+yxi5RfTZ3IQg71rcNepXQi5eQ8qQ4tkMbREzWtu
LZSNTADEppguORpvrHULOfJmFSm9g0/Z5LA6QkrV1SWu/ip9V++vlDaQwL7h58r62C4yGnMxAf65
ibCVyce7QbSe5Fr5rmjxj4wc1KeMej18p8Z3FJwEeopUOPOTawKmr9PjEXpQ9O099BBBPk/9zMDA
a4BFdrv2DiXIF0YJSPA+eA3lg4H5OxNef2MlwxrEvBp68mDJgdCHe7xHclsyuwJRUna1PFp7xUU3
fxWKHFzHdiq5cBUHBPPjYAQkCFuZ7ZkIiQCmE+NGQrSx5UkzyLVwEvLImisdfLMGGEzbrGUWSpqg
Xk4pgl/JsPjHRtuCINC60oybwKGLdsSam4XYgmu2h9crTjr5obWPKmjaYm/Oxd3IL99EdfZIHT4x
9wZiAaNbLjxeIJNmcJ34faO1loRvcbyBP2z9PPqV+u0nY6Ct0Clz29DDv24gB0uegNw83J5d/rgv
whkc+LRhR08XUQ9MdH3IANGHNzTENzH0H2SWDnaxks8etN4XbjKiHF1SUJG7OlLISxDnlMttRgQz
H80ikn9c1qKfjSIczu1EobxRY03/qPEEamrObcZn7Z1swrPziM1yjYnZqyhifkqKdsZUgOzzlePD
SE2JQKxdrcqtZqFubJbf9n42Kla3NacQDqyn5N5RvGkhQ5Mct03AkHW6hDagbl3xHSoxvfcEmArk
0YkirCPnyGohNmpR2Z9Uwt5v87v6iTCik7hS0XKtUouFFqKHQMxaXU8xcpJ5K0BloFKpPECkodti
Y3b1JiWR1YYONF2zcxwCvheWWHyJOPV4cGlYF5DYG5hwCbrr0jwydBxupxrt0JhK72usVBHR2BZR
Rz2V3aqSCfcvV0W6z5Yy/TwC09AOS5gt5h+dF3uK48sSy8LXiF08Dt2Crm2J+cWg7K9Y28+7zzk8
tJfxXXue8QihBJccOA+dipjLl+WlTfsJAjfaVV3WZNYhgL1++iiM2AiI+CQh8m5Pc+pHh6/KBr6I
EqZeNQxW+6oZ9a7tiLQLVw4BjhixBL9MGIKlp52ZPcsgTDj/+one1DpYchy6HdmvWS0rwU8S13SU
oT9Uf+IAxazB8XDqanJYBADXmXQoIEgPKVg8eahZsWvL/CKCFyikK13Nc7eGEw3ftppo2KPK3KBR
pvVJRrOQIc+PkYZ1AkSIDmNAdTD3x9QGjbCjYcu3mgIdJDDjyUOdUWovvF1LQ4zkvPCEOJ+U6nXT
Lrm8WhNluxZ4GyDnmONt3Smk/z0CpZtgRLQx9S70dD2C983v5nk3IRElEC2zywdywLq0sjdCKRkE
Is5V5k2cni3vZjWfEGm28osFPDZYQpUm5cLiFjNPn6lGeiwn/HBr7S0NALjQ4OVzGaYw6Rb++JcP
cBP5VZFJc1KGaK6N2hkZwA+cgSKnHTvuoQLiG03rribH3tEb8Qdqcpk5HewStjzFJMrcDQrYHUTk
sw+J+SV1DYw2nuDO12LoQAHJq4/wQpipj2vWesEZ9byOUPjg+qyS62GX0YpPUqouvCRhAIB2ADr4
TvFh5+nAIE6hiQk10cksDl4GUgYDpDHLnfHT1U0kE8TjILkOfzPc/02W85cU982tLrPBjWhDMEwu
HnxuKmQgJuKc224jtBEZ6xCuEYrZpOc9atobbuqjLqTOSmF8167NiO0aOOhOgTOOtKAbcvpLYRMO
1zxY+GTiHJrR/SxmG1fEfhLs6S7HB4QCURAtpJzx130V9rFV6uiz4ivNsW5DH1AQXUEdiidjrcLr
KwU+C2fKWAsofocuaBHgkLPDVYVFiQWxXqkV00uZSiY6aImOOBVV0ptcsGe128K+phRic/QgQlaF
0kFF6zlXbtKmGL5JN2jyeY1q+LXEBUc3EAnW802YzoOp3OldaGg7BG4QPpDo0aVmhaL26/ulvZnC
xJ9jGRSdA20t24rZRqnjCI+9QPULGIUniyLAKH8iqM5rUdIlP3NcH1cb0KCELx+tk7QbSnodgRyi
yOnL5KfGgoZa7eTFM4azLN9m0Ht3mrvE9aZOqu6N1pD0SuCqogBaSZD61TLeJg76JAAJ4ZYdvcQR
suOGzcFZ1q74pODgHqqHEfishdoFT5im06mco//GhZOEPedmms/LHIdgEuYq5SDX5lZbnqGM3/Tw
q79NMoLFex3YYhlM7WszTZ2NuqL9MUOdF5NXwkyVu6z4Jsjpb+PHwUcsrA+lzbOq/KJb/EtqmxPO
dFQqqUXIp/vtbDzHYSnY5W1R8pSMECiP7sb5kGRYjOhOvXF7P00efiqO7fNIVOI+EO06QFO5inQy
zanUJmg0WPUjg11i+lww0kwFNGFnf8JZF7Bivi87PEVpqfv//6S7FcA2fZZxTrFdJiIlH/cEg5q2
H7dMrJHXPOXFPiSBWeeIo+44hStGjEXg911MZoZL1oYAtkjgHWHr3QSWfBcQ3/QUI1Az/Finy8dk
mJVzdRNNVbHMqKCIYDkFyabCKS9XWcgcSysLloYfU9gyr+cv12AwQA2PAs82tut3nzdK9/Z0lADn
CfoMGelx6mipgH65bpMV1wYmD8GnntjPSkGtrUWJ8chuLPyf+Pn8q0QXFV5Eb8JbvfYpLpCbDshO
TBLJ8/2ccaz4jvPBVfuxXDgfHMNGR3oulPFLT9vB23jh8RmPl/IwXmcb6WZOEm0lwDsM4H9n1NHT
Y41qj0SwZOro8DNH8OsY73jlHGh2AAG1AI/ivj6wkdA2TieWLU+ccCBZ5ra+dkexrH6pYAEFw3Xj
ynGYljPbtxjPGtm4y1DnU9jGR7XRoE2z5bo9Q4Brnc0aHrv/jykIAt9xW7jKILE/Y0q4QMc12838
AMMOZhWhbu2JAKdaKdj39mP0xUZ69TRze93ivaAnXeqfUJYt9kiJZcL+LS4necAfXmNTB57on7lw
wFTjJePkSBweuWCtg+Vd9+LuenmKjXi9NshI645Bn6F9Nt49G/lSrVMeLNxNnkjs7RGXa6/G8F6u
N08CCLNf/qC6co76pcOW5omfT9VcLmva0wnz5qNg+VwPAMrRsHJlEGT7KhzbqpQ4y+/LEJGKergt
+Oa3U4aKyA3TkbBh9p6meoqUu6qFigFN/4SHXr+N4vRanUFGXVaCIs9wpSBactkcUgzAToHGZCMO
Mq9cww8xpwCuu1VDF33l65xZPc4xcFVDAfFsfMrhiD8aziAfBl2GDCQuR31p3uOyaLKSxevsmCGs
n2XhFIZoOLAhohgxnMVUsEM55BtbGsT3Oz/4jjB+MwOwKzPrQTvjOF1E1xD1z24YZw+Po0/rvy6T
5TPxQwNLx64xdoPrvSwQg9DOIj/FeOJHJsgFh5nhgE+8yS925+mT/fBw0i3lqTxJ9Z+OohQCd6RW
kdekE6XG4a+C77wzJJSrw270Su9iJJiu+QS+FWwGlX6++EQh2j1L9q9N/j28QQdojfmBRtL6hSTL
dWJpHIgeWm3gGuS4r2K6qtkJFKLQNOyYnW2Nu/RuZ6VElhlFl685s2ic1kzDps60i540CeGbMmSi
PRlpDH7JfeiDRHWEHAQKxpw8fhwgw8OoRDhssSw9SHomv4A+XrnC/Lot2XiT/29Cyjsb1a1OLECa
L1o0VbnHwSDxRYzsT4WMm1pKMBve70P3utVGwPEWyl45jnvd+9iUNaq9pDbczzBPFbWwUHtnddin
Qr2LPAudg7DvuWuRCAXUL2+esEhpUCpxBeYE4XWRAJo4JAS/57Uuy448f5qdySh0VfeER1uL7Hu2
sTwmwJiIDdfX5iPtdWEForAAXCgQuX0Q23rerX9C/Z8f+rgtUxh2NIlnImyO17v3zQAZuCI0y6bD
Q7vpVc28qq6zraKa8YGBICYbQVe4eXWkEc4DcljTBBgGLpXXljTcSeFeiSOkveZVd89sCBa0FgEV
o+L+GKKOe+lW5YDQ3I9Yf0FC+0CDuylZ50ryVrEDcDn97K/ulC4nLsinSA2uVqr6D3j0MW97Q2Vb
forZA2HLNMRX3SfIEEOtyTvWiPd69zdpFcrQv4Hvi4d20sHe6TJW8HXzz2thyXQ959T0Ba4U60dg
JAhy3myKi8ZebYVIioD53SFlb5z8+7K6Qw1aVs7PWktrlCF1OQUrp6d/ETNT3BghECtyw+tq+erj
yGP37RtMuTkMAvdaGpktHzcvZEwtm3bBenR4Mtwv6juVgV/bS1qRpriRbWsHuI8tBHXZz/j4X8bv
BXKYygtSDwdJc5TVl0ozvrL9eBUgMSJeKtGui8fXz/Q+bXr6JgMeIdTR01jninvtOPpuXAmTWieT
hwKzjW6e2J2GksXDH4d1e2uekW16yH4n5YhhZ8Ms37q17oylM2DnGvjfFmAPv6QUIjPx29G2KtgX
rxB/g9kn91tU+OgCIWd7KPT02skRMjd02D+sJIHThvEQUiyauWYKKFNIHW0hG4qHCbklz3uW5N9F
5izcMbER2qCfc4mLxNJc4q1fui6V26PaefkUu+WVW4FnVdrMQwgTBvCycZg6uEBhisblYhmyK7Tm
u/HO38P7Jd3W6S9nm/73OQJ+IWIe2/xzNO9/FXDTgVEpV2OMJbztF5JhDYaXGFBTVMxt2SM+gutc
LZTqM8LeRODvAbXDXfcgdnoXGp5qbR9UO8CclEYQS7/GgqqCGGDhR9kCjz7TI0uqGm8ERL0OTEbM
wt9zG+SPM75WugINNw4o4RL6MghwKdCJn6a+5zjWsnLfrmvJt+IIGxQzwbv/CTv82DLddm3L3yCA
HUSlCzJt/1V+iZc3OdQDOqHpyEd/JGjv0xrNs3ZJWYw1b6Y3/hwCzoxUZV6aCFVnwgT1KUpkWND8
tisB2ee/XrzG40A3g2Ji+CNuFSqxrMOlofkEUnIlfcA+VWbJVLnlTv1lfVWY1K0sOZLXYPWUhrX1
FIHElwrTkcGheiraN9bfuhv2IdVtIs7+6Qb0/NTR3sAKUxMjCBNIMkDcMirUycBulLms+VVld5/J
bU9A6h6p49RdS2+8aoP+rMjN9VwnvMG2RB5o4NGUfk2wBOq/18Jcp6fbkiJQaY6FzH31IWnxCRq7
K64oXXldlyml8YnzJWwMRqL1styZBIowIt5c43emP8UshgyB/pD4pVBCyyoEONT9qU8jNzMeKtt7
9F6aEKGeEv2ZKvPv/BkiGUGupoTzWyy5QrmI2TnhoQp1NL0bQ+PRWGDxlokl5uF+VOAJbeQvVg+j
CJfNTHilus+66zHwrrw7lOdZ2Fj9j2cOpv+76suCgPNIWqmClQTJglBi0ZdF7BUQEI0kApGWqhwr
FgjJGGjfQl8zxvha6QbjwO3NWHsM/mhzoj+10zEMcnybNzpMvoBq/AJPYgyO0Vk2KUXe82JnshZR
5zAxSM5EKAIurpKh05dIe6LpOqC/D9IJ/VDdVlqIgTu9Q5fctZPhySq467ZAE20Tc276amfMQj8e
AIt8AzILolitCQWtErvD7+p069ANjt+6m1ZRRncWcLoNQSVDFcE9cJ87rLVp0v9t+QfWXC/TA/Eo
z5UfIqKaMFjvDTREX8mSAZB6Hx9gtuNGw4etV+V4VYZqYzVKpxnKMOT5uU3Q5FOM4kH3afu9WlOe
Djb7eCb3XITpgfYj4TRKl/h3Ys91thOdcgQf2rcJa4VlqmHYGReB18D3ua3IVq5o89dk3S28W5a2
lH3y1bRtgVBlbliYNQx7bXuFpLZYSFVcw1zY8k6BCKuuX6IwcUcC79hXH1ysrMFOVZyoTnKHjZeD
KWMXn4otPK+XM76LLGVw1X0m6CulefMIT/LFVw0649CPj8i1z7c1EqqZTRm8xM3KE243ygPnKlkO
aOrfSj1RGtLQLbjBQkb2F+qQP3vjV5R24q36upG4VLkG5q/I0QYhv+5znTiYSgd2evhUjZSCfbIa
wjjh/hUyZkpGVpBUDoSSTG7/UXmoWVBb3lWdTZ4Bf7rq+uDutJFk1N0hGSSr3wvOLY5qzTr4vVQe
Qo0jS4i2nXlI6TyqJqeT05638elfKGP0IMSId7Tre+8ucwAicr65coK5dSssa/h06YDPzATDd8Z5
ybK/pA5wdpWX9m5XoXIZQ6ebUnm5g+7/JBdZDkd6/gKns20VksfOuuhJf9FQ8NbCzwcqVsUEXMCh
c6rMDRpSxHziXiaKmWo13ZWjjmMsliuwkh2NQKUGrsT5tqSJkk+4ZjLjg88W6W+ZDe76iAieJfbw
lg6D7xfOynuEFu+SVKjykaZWtDcZ1YCsuogJyV0EF81xRn6ItDWQqvP6lqtM2QPkc4hJAEcDEesG
Qvq+K74gS1xwzr1BBGNvZX2MVeopDSiTskuxDfRzmawUlcHMz7ye/+9y14IewFfgG8ro7JTMMjgD
2am1UZhCW6D9nJ0wMnHFWXYHD6+F+G6ZQ3C6cAlZmIfdwTLaRbG8eduvwUbMzS67ZkaGd3FbcoKN
lsTaJn/tIpPZJ17dBh2imHdAqAhECZcBA4xmiwdmgnR7XHOufDtB8Eu1fRMVm3NhX2MZMi5/hh+a
oVX56RCtkkMQ0uDhQYOZq4HHCqLFE6/jAw9lM3COqLcLrKK9gmaxSLCwifJu2xL2fXHDwT3qbbOv
zuofADuPS21IYX8Y019GJ8sdtX0tSYBdKDzOAWL9tT/F1nd8R04NGjyQNJ7uruzLOopbHeNQcSHN
N8TBWfoYqY0JyqBZSDL63+D0LIK21nzFYJd34DOJYsL3mp1BbkbibjA5VVM2PgjZpdlGexxHLC+8
GUzkhdUXmj1xRmw/g4KFBY73yS9M6YO3KdheKDHi8WVozOxM4ZOriCWCmODrOWjmDNI4a2YgpoqQ
60UAldQTx3IIwoSJANNje6CJ9FKYpHRCFH3DdXok9mBBMQg0LKiNBTqz4/8Fi7WGAXqx1bwjao8y
zzpxQOQKJFuioahGRIXJw9Qpy+5rTzLGqyyAxE5BoNwnh3DgMEm+PPtIhdTe8uU+zLewEN/5FZta
HPTysyjYg4Y/HxoufXbXm9bTzRjE27eGwJ+Sp4x8NvmQzjY+wn2URyBYR919rpPW6YddYO2Pvh+r
wK6ODt9BvD/Hnqr+f/GJsd+i5MIZ7m8/IJtGCIDjWfSv3Tv5iUoJVN2hASgShLa5khzvuZ+QvuU4
/8bjznoEMQvDb4Onzc/gmvnkuI0RbdfKVkvW2O1FfBjT7OUd+BR/HZexCa/wipfiLutP7YpIn7le
L6BYgE9UkRK9p4brCoVXr5oKXdXRcq2WanVhcVk2m1gawJ4JMEOlXILJZWwKr6NtHBH2b3oIqa7t
WfYAX6JPNRp2b/2RehqBuzQd1PdBcATfpv7b/FrZ19yFd5mbzDXwPFp9eQjfXHj0iycqE9WXga7d
5DG+uupoECxZtMc7IX3gKw0pXYkCLSUr1bNb1qk2mlS+Nk+OIFlVtMcXe7FEFXv5DWG4uXMKM+hy
trehBt1wOGBQuOltW0c0EP7K99Ll8jo8gvuWlyEzc7JwmX09mqS/ajxQpudDbLFwsbF2WmqM635O
QXGfUYleSadGjqUq2gG4R+wYnJCqKa2KHRP3PyXG9kzy7KZmayjcV4zbmPmXwRZJHhecpPwUWYQY
/T2yzX0F40Plmq+JRgdKGlIHQmDIzOmUbrcYQbe7WsM2ewbBemeCVT/K1tBWbeLOl8v0fVAYFzNV
1n+2X+eSwbRGMpljhg9nXAcF5VLDn5rn2fkw0GCjoJFY5Y9TlW0X7vQVm9N7xE0VvJ204+we3tE6
DN/a683LC0DrmmSqKbwp5U/n/Wg4IHqipiOBI3lXSlYRaWNsp3+8+/bgMLl/kseiLlU/VTX4Ugcr
wx0q5ha4/rqCEIYM5J1OjlZPa39QDhb3opxrITDy51Q7S0MhzDlo3zF6Ei59fK0M0kTwmPIjsQF8
P5sod4BmR+bEnAl1wMs0SnRgQSdB3puxz8uq6img5JoBNvEEjuNRa8C9UvMUb/oamK8UrqQ9r+/n
aEAmYptihcTlsoIPfD23jp/xamdSjPCVmrDmxC8M/0T0DKLahqoxWiExKQh8zJqiZiwBoQXS85Xw
JaWUfBEgyfnh6I1FVOXK1awYV8bn171LwYnBupkSM4Z70um1IDHGiZEGKkApOQxUMWKH/jOSC6E/
uXn+FGHG51sjBIJ92P/mOM0cEp9u53n0FPwaR9TEWnHY4ZFHfwl3kWNrCb2tlLzs2PLCPVE9VMld
K9w6lR8zJm96xMa1ArXKbXwOt9UHPDqq9Hzg/kelU7wFNuGgECFNM2VtM9OganQizQsICRnsshTq
0erqexVXp2Zu1pXS5JaQ3BLDqV3RzfKyabdIzQiElTjEhnLg5uP3cm10CzKTC9slTxlxLydqVY4g
vuFDRCGaJXHbqbq8XkOdQr+eub6lu0ztlDqElw0RoV3AqZPLBncdqvCuPKSCDnmULh06JGrJ+YSY
sDl3Zq3n0fYouXnZ+ogZ9A2wv4SQWYPBmZpO9045fA8yIHP1ZH75h2+5bt9RCjsJfI2/vZtetak6
zavVyEYKBrD0ovcaiPDWF4y+zB2qfJNJwfOWOmDKoZJu9+crUwUo2ZD6CplOZU7xfN4R4InoYc71
SHX49DOe4hxR2h20EqMv8Roe3rc+tMkZe6ESTgEo2sWlZshcMNJoQkuJ0A76kixDPUjohmDszcwd
R9GLEqrrIiycCUpqm9vjSIIuVu+VIOLkz+1LEmbSSrzGI+sDF21tiS5ZaoKP4f71XiEvhpLlA92n
YkY400sKtXrXDkzDLnd1FIQ7T1Xt84nDfrKtoMQfq0CPvqxn+70TlMyHH4Of4Okk7O/7ulS/Fkgv
kqLDzH9aFo70AX1a9Idrjr+jvgp3ncjd7ItZhnp7xycQyqI4XgYXvBKElOCxjXsHFjoPpOR62jFe
wFmL4JEB0eYO/ghsulYLwiuGYjd7YqSVbWWoEm8/Hu2Oy4XFn1/DaeAoUXC/uJh0F9oV0cs1VbRL
FUV5N//r9jybSI4j7NdiIU7P7tWBn8BI5MnPImOGPxtbu6Cx/LL8YhmG7QbCVZji3WJ2Ke4lI3T6
Q+v9PYUYyoSNIyxxYb8xM2F/yRmmOiWt08oS5jz1z/XT2ZB7DZF/Np0EvG864hwBLV+frKU2YKHH
QUtZVbC5fulpFHPTtkK0bPYh0uLIeC7sLtHiRSUe8RpCISN7H0Q66lAYMuiyodY6kWDEVBoFwTkO
mRozyK4NF4MEOrNp/hEstmFc6FkQo8WQbwmiFKiu8/sWVYCNDD9X+gty+7HDKkFcsiH/Fh37hOmD
gcRSSv3Ga3NrbStDACQ+KILMk8B9dUGeU5lD4ISKOfYrp1QvTWdp3bifnZcFqUryLkJZ1CSD1XNO
dz9mgbemX4TK+ik3ebFL9W54pAI0NFDnLLxfGCjhZZNaDihsjwtvftfNwEhWhX9nMbrdzwUwHDVL
Ucxprj/klQFtxgkxpjGn1cX8bWrc0sIX4oYt9as4bq9a59YGiPQxdpBL0EvBRzuPsxlp9GLieg0H
CkOc74Wy3FxM6NHuxS7KzVv9HLxLpjXl28jMCqHHtGy/DoMO32qn4WwoDqatV1RzjpOhZtix3T7K
QRy53H7hUYAiZbSlG7SmUuUl/135zM3xcjy5NAVfwjrLlL48mHNq4U7KVbWd+XByiLxem3RrqZR0
QuF0JNNUzAcZ0WvKZ7Y0LADTYeHHfNt8UoInDx15r/gqLEd6VuYH/VH4I1rVUyWg+u7XGC2q8zfQ
yFYOFYjID/7hMNR7mgm3RfO7yhL6f/Z0LkId+gSnzm8KR1JDbfFM77WVNCRQiFBOWyYaT1u8G0UY
9VauMPPxFfaS1FguzDAQgAeBVThz21pL76/3N/J48HKFuCi1IHfYcOKKdLWCfm95j820HZJv9XMD
SLK9P67Lws/8fa01ZDBA/LrZG0/ifRfYO/CGz1Ob6c91k7Wzz0Q0QeC+/1G289mFuKgMPKuGhMO/
qurMicikIwHNZmZo3b44saky0WaC6ejm6GxE6Y/Fqvdnk6fCKkbEjqlTphYWVduUeRIUBQrun4gu
BD5ct/Kdc+qwn3GJu7znZ1zyQaZiYG5BBX/O+xGovq0vdI5ZnNCdKQSXEWzDN/FdMSkY/ptcEJd0
ia6jej4JkfPMiWtgZSxEFCnhNoaRcHXK4Z+XP69IVLyjVk7Fu87D26G69Y3IoVThdWdWE2Zjnp5E
UiYjGn235LGDxqBmkS78tHTb3A1ppua58pAdX5gxUgm2VI+HpMwE1TResoJK4vX+Ld6HtHVrKjxu
jY2v1pkC76rGSg74geIFVAOaPSzrXWHqoz03OkVrUmikUgm98S0uOxN9eXMetsFA1sPkQEhCZoLS
9KMgDDbWAcGQkLnlwqOJ42lRHz9qU/j4yBSUkWmVDQtK+I5WuIQP58DQvotQPOnWE7afDn3VMu10
qbWbJ2SYL5kX2KEgz9eEjCKUOSWKgioT35ghO7faQzrBxF7Uia7bLa0+aeAgPlUSAJ9DJVzzteqv
HqvM59lVUtKnKFXBQKN/bLUNvkXAVNjeflfpKN2PF8j/4M4W5n0PVJwXYSbw1+g7zCM8iMykkDrS
Hvr4gDYKnmzt+oQIDaV6HI0pYYX6Zv0yf++/g42zv2qu5b2MGmzsDyMCGU8VmZa7Rfh2PqH3gF+Q
zjP7aJKobHThqnEPbdGn9l7EsAWX8YcyjYDy83COWskKSuDoz3y6uH0A7XMoD+oSrdyIeGgC2yg+
X0Ijt/pRwv1OzhzYIIWZAqVyfh/4gEwPackvULoU1yOPTN7XCxBQmaWNN7boCphoIQ9jUxEkacjx
PkOrfsJpkSn39i2kYx2qC5fVXRmd/Z+WIpHnu50cWBE9EYUYY9a2vgMFUU4is6+b2jyeSCTUV0BG
l/BlwlD0IAtI4Nd+NjV8DKcA/C/1zFigVgh+KzAbfa8hXacfA10RK128CWShOv91ZIiMWceFq1hG
p7WjGGXLJloYUo78UgHoJgXEv4/Osk/mRPRyCRHBXD4+hS09oFrHzT74fg+CIbHHU8f3O8JAmZGh
8DG8qiBvUMNvrhmE2Qm4plUSr4GwTPAeH1h9jjdAMDuJbWg88VYurXpOtjDl67JIgP1+tySPX9YX
VaUD9p/RsguJ8hoUNUt22RPTCrEIESAr8QISGIE/+QzmyLKZptEcg2qRBvGAHQKQV5X0J0m/VJZ6
+tnNa7Zm2+9OeZIOsTbjDiT6gqSssM86ZW/gpsREGrjfJLbyvaqrEoHu3eBKwhyiz/mZpco0JGDc
VHsA7ztt/QLw8mdh4DQIWAjzWNTJekxROYkdeJRmDn3HSuTDFeaPwwof7UJ7jaVx/eMd081656lf
u/fU+FxBdrs3q0vR+LEhx7vE4KIW+y4h0sFbwkUrop/uzXmZyDu15vslsTLZoodpw+1csKsD/ML+
NiHvq5VcX3S90Ha3OxkxAfRwNnI39NF0v2Dsm8zm65Wjha0oahJzGLWEubC8cNQAdRNxQm+o3Ehr
Xu9avkWTksg8FBQMgNlor50949F2PRqCEMLJRW4Azl2T1UdBw/NZr0dkM7K8u5+4yX1R0ogdX6Cz
LSdFXbf6wRWJiPEt+x0nt10r4j6gRXYhiFs/Ct00K2Vma9s1REQBtCcE28ttOmBfLvAhFeAgAD78
9E/SAD4MdUkeC8cGdk+3bF8pc3SYFRtEQ/4/FluY0JsLTQ9WeXEwJi/gkweTER0AzyUUJe/xY0wS
Sfzo2BbSx2HCf2ahLPrl7Lfzb8JYtNpxGHIQrzQ1vI+lCGlSg/L6HuePP7eCbJS90hxCHfe0HE8i
P38YY5tnlm7zPpz3McA/eF+yDHb3b0qK/SuMI1ZsoJcFzzUsuKU0AGGyU4a4D2CNe0Buzei/8cmk
uqCdzSonQRbIsP4w/BuMm5RFHg6PJ1ISZPh/uyN/hlrIZ24FZCOc3OhhnmNXwzd2aNOOiZ264yXb
vJ9y2V0qyEaicmai75iM5qC0SdHOpf+tRANbAdN1mvcuQf3d54xpzVYpbvpNwnTNCs7r04NYYPqE
HnNRsmpbwFHU4GbdJR17Owqx6NTMhhvSIUO4OinOOhX0vY4SaOb10RFtwwpJJpS5iIcNg0eIhuab
vQVQ1HHVd3sFrnKfW87hxOTZpcYVWje9zGy3utMDjGyb3Zh7kqI0nrfUU+7K3BMxi7oQTqaBQeeJ
lRQCbGftzlqphbj8HA/nzLEUHuNZNH0d6+wGmaw9Ev/r9i7P8kSGMG7QYlEGKTPOg8+JAnUgFe1D
ivsEN5JTHGQsyZoSu9pRfq2Ta4v68Lu5fIIwrlLj5KWLtd1xUAxuiHNb3YOMZe2Digx2yqfajWhF
pszzOcAtyoL5LPf4WjTFGWByat+3rpf/vFFZ8XyCSxjpIv0hapHnR2vLrlF+VE/cveCM7AwwlMHX
OaBOV94XPJbHaSaBXNfpY44APmTxRL+W5k0GKmCSqFiC8Z97z222vlPZHWdfej7tlBXIK3jZz4iQ
U3vJHWNxImR10llLRvgp1fNtNmJKlid3BTtJnJrV4l/S2gJ6qgUSnqMioG/qTkEoofrJLjG4Eda9
PP44T7RTd82xKWMTy4sPfTyDWkJ7fPP0TICpofxnjtNZodZuSZHw9JsPPWyRD3jdpw0sR0/Kayrl
U3PNz4mpyPS+r9jJulkojSBZVP1ts8PpheOetIQMbZGsMT9w5Ocw3A7eD3OXNNC/kkvgieymdMgS
vl3Te05h+B5Q5zZvorV/prm2suEXZkAojv6zrhyetVATeq6cgTfkZUeZHbJaz1FZWqwhHMQZm2ii
qEAAfAr+jsfx1ursFANkjOs7/LE8zDHS8TNr5pw/s6PtDWF11fHxZ/LpvUG1axsHX/faUrqFW9bC
kzH7diPkl7CpqoqqbWl7IgstFDyf/wVjYeju7TFGMtEZSBwFVcwY+9zPJimm3M4Z/D46uEjwwSB4
jJSh7svcoEtwtxZcvKmekAuVCKsNYMMXDhq0wWiJJj8AIblXbXz7n/RLEoYkcDHAK1iLJlRrqQpw
S18TMNh4S3u9j+SEPUTAoCh/Fw0LkjoJjmOdywIkZwAEsqbjPAwgKu7z4ReAmm8cjPlc36DnVkVU
GYqS0gO2zYXTu+M6b17UFoti6RM+1Sl0AYg0NUxQXTRQP5nuzcFhS7h1nNFoDGWY6dXsEfjUqcvT
suYF1WMo88j67KawNpVOQYcFikgADaP4kY87n34iBxuCPZrKNRjuaoZEwq43IVhT/c/grkgKE51H
AVJsDm/M8l4LvFjLfMX116VGJxaS5WQKABctO6aMlvDMrxcmT4jFnmwmy1cEp8sj66fiS+Ydd9gi
s7BaXA8W4gbKbHyPrthCxsO3rwIoAawpxrMf/ly4o3gi6zL74T4isGCqc60HPUsW6MjgfgDbiMV1
pcGHzH1SSdi7UhaJ3fYlHK3OflNu4H9YBkxp2/7wXhQAk4IVvwn/RRnvwTvZY2eXEcMi7vDGXyKG
gsj1JNH7N3Qt1G8KfTX+KGKvt+HXQ8Puk3HKlEAD/dqG1v2M4HqmpOgxp/4yQHnwL/c13DROApUe
OxRaitUTwv48t948IVII+ZmBrV7Cw2tRKl5a5t3YDPQ/iZzYLC5rJTL7Lt9TOOZPQiVqsJkWdz+L
h+XzeeRfnu4SnY0wyRElxrlzs+MuI3O8b3M8GC+U5VS1uTA17c+HrGiVxkfHrp8zZuEe3Zr+8QfF
9KYN+NXREtSXF1scT4YUzvqffO+WHU5ktzyhWskkypvFkJAf+JxoEfJwl5yAXxaL9CgIJINYLuFH
ljIrToESclD2pCEWJEi6jrfQOA3ZV0o2EUWM5Q==
`protect end_protected
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library gw2a;
use gw2a.components.all;

entity WatchEventsCore is
port(
  Data :  in std_logic_vector(71 downto 0);
  Clk :  in std_logic;
  WrEn :  in std_logic;
  RdEn :  in std_logic;
  Reset :  in std_logic;
  Q :  out std_logic_vector(71 downto 0);
  Empty :  out std_logic;
  Full :  out std_logic);
end WatchEventsCore;
architecture beh of WatchEventsCore is
  signal GND_0 : std_logic ;
  signal VCC_0 : std_logic ;
  signal NN : std_logic;
component \~fifo_sc_hs.WatchEventsCore\
port(
  Clk: in std_logic;
  Reset: in std_logic;
  GND_0: in std_logic;
  VCC_0: in std_logic;
  WrEn: in std_logic;
  RdEn: in std_logic;
  Data : in std_logic_vector(71 downto 0);
  Empty: out std_logic;
  Full: out std_logic;
  Q : out std_logic_vector(71 downto 0));
end component;
begin
GND_s0: GND
port map (
  G => GND_0);
VCC_s0: VCC
port map (
  V => VCC_0);
GSR_0: GSR
port map (
  GSRI => VCC_0);
fifo_sc_hs_inst: \~fifo_sc_hs.WatchEventsCore\
port map(
  Clk => Clk,
  Reset => Reset,
  GND_0 => GND_0,
  VCC_0 => VCC_0,
  WrEn => WrEn,
  RdEn => RdEn,
  Data(71 downto 0) => Data(71 downto 0),
  Empty => NN,
  Full => Full,
  Q(71 downto 0) => Q(71 downto 0));
  Empty <= NN;
end beh;

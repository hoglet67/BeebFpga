library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity saa5050_rom is
    Port (
        address : in  std_logic_vector(11 downto 0);
        clock  : in  std_logic;
        q : out std_logic_vector(7 downto 0)
        );
end;

architecture RTL of saa5050_rom is

    signal rom_addr : std_logic_vector(11 downto 0);

begin

    p_addr : process(address)
    begin
        rom_addr              <= (others => '0');
        rom_addr(11 downto 0) <= address;
    end process;

    p_rom : process
    begin
        wait until rising_edge(clock);
        q <= (others => '0');
        case rom_addr is
            when x"000" => q <= x"00";
            when x"001" => q <= x"00";
            when x"002" => q <= x"00";
            when x"003" => q <= x"00";
            when x"004" => q <= x"00";
            when x"005" => q <= x"00";
            when x"006" => q <= x"00";
            when x"007" => q <= x"00";
            when x"008" => q <= x"00";
            when x"009" => q <= x"00";
            when x"00A" => q <= x"00";
            when x"00B" => q <= x"00";
            when x"00C" => q <= x"00";
            when x"00D" => q <= x"00";
            when x"00E" => q <= x"00";
            when x"00F" => q <= x"00";
            when x"010" => q <= x"00";
            when x"011" => q <= x"00";
            when x"012" => q <= x"00";
            when x"013" => q <= x"00";
            when x"014" => q <= x"00";
            when x"015" => q <= x"00";
            when x"016" => q <= x"00";
            when x"017" => q <= x"00";
            when x"018" => q <= x"00";
            when x"019" => q <= x"00";
            when x"01A" => q <= x"00";
            when x"01B" => q <= x"00";
            when x"01C" => q <= x"00";
            when x"01D" => q <= x"00";
            when x"01E" => q <= x"00";
            when x"01F" => q <= x"00";
            when x"020" => q <= x"00";
            when x"021" => q <= x"00";
            when x"022" => q <= x"00";
            when x"023" => q <= x"00";
            when x"024" => q <= x"00";
            when x"025" => q <= x"00";
            when x"026" => q <= x"00";
            when x"027" => q <= x"00";
            when x"028" => q <= x"00";
            when x"029" => q <= x"00";
            when x"02A" => q <= x"00";
            when x"02B" => q <= x"00";
            when x"02C" => q <= x"00";
            when x"02D" => q <= x"00";
            when x"02E" => q <= x"00";
            when x"02F" => q <= x"00";
            when x"030" => q <= x"00";
            when x"031" => q <= x"00";
            when x"032" => q <= x"00";
            when x"033" => q <= x"00";
            when x"034" => q <= x"00";
            when x"035" => q <= x"00";
            when x"036" => q <= x"00";
            when x"037" => q <= x"00";
            when x"038" => q <= x"00";
            when x"039" => q <= x"00";
            when x"03A" => q <= x"00";
            when x"03B" => q <= x"00";
            when x"03C" => q <= x"00";
            when x"03D" => q <= x"00";
            when x"03E" => q <= x"00";
            when x"03F" => q <= x"00";
            when x"040" => q <= x"00";
            when x"041" => q <= x"00";
            when x"042" => q <= x"00";
            when x"043" => q <= x"00";
            when x"044" => q <= x"00";
            when x"045" => q <= x"00";
            when x"046" => q <= x"00";
            when x"047" => q <= x"00";
            when x"048" => q <= x"00";
            when x"049" => q <= x"00";
            when x"04A" => q <= x"00";
            when x"04B" => q <= x"00";
            when x"04C" => q <= x"00";
            when x"04D" => q <= x"00";
            when x"04E" => q <= x"00";
            when x"04F" => q <= x"00";
            when x"050" => q <= x"00";
            when x"051" => q <= x"00";
            when x"052" => q <= x"00";
            when x"053" => q <= x"00";
            when x"054" => q <= x"00";
            when x"055" => q <= x"00";
            when x"056" => q <= x"00";
            when x"057" => q <= x"00";
            when x"058" => q <= x"00";
            when x"059" => q <= x"00";
            when x"05A" => q <= x"00";
            when x"05B" => q <= x"00";
            when x"05C" => q <= x"00";
            when x"05D" => q <= x"00";
            when x"05E" => q <= x"00";
            when x"05F" => q <= x"00";
            when x"060" => q <= x"00";
            when x"061" => q <= x"00";
            when x"062" => q <= x"00";
            when x"063" => q <= x"00";
            when x"064" => q <= x"00";
            when x"065" => q <= x"00";
            when x"066" => q <= x"00";
            when x"067" => q <= x"00";
            when x"068" => q <= x"00";
            when x"069" => q <= x"00";
            when x"06A" => q <= x"00";
            when x"06B" => q <= x"00";
            when x"06C" => q <= x"00";
            when x"06D" => q <= x"00";
            when x"06E" => q <= x"00";
            when x"06F" => q <= x"00";
            when x"070" => q <= x"00";
            when x"071" => q <= x"00";
            when x"072" => q <= x"00";
            when x"073" => q <= x"00";
            when x"074" => q <= x"00";
            when x"075" => q <= x"00";
            when x"076" => q <= x"00";
            when x"077" => q <= x"00";
            when x"078" => q <= x"00";
            when x"079" => q <= x"00";
            when x"07A" => q <= x"00";
            when x"07B" => q <= x"00";
            when x"07C" => q <= x"00";
            when x"07D" => q <= x"00";
            when x"07E" => q <= x"00";
            when x"07F" => q <= x"00";
            when x"080" => q <= x"00";
            when x"081" => q <= x"00";
            when x"082" => q <= x"00";
            when x"083" => q <= x"00";
            when x"084" => q <= x"00";
            when x"085" => q <= x"00";
            when x"086" => q <= x"00";
            when x"087" => q <= x"00";
            when x"088" => q <= x"00";
            when x"089" => q <= x"00";
            when x"08A" => q <= x"00";
            when x"08B" => q <= x"00";
            when x"08C" => q <= x"00";
            when x"08D" => q <= x"00";
            when x"08E" => q <= x"00";
            when x"08F" => q <= x"00";
            when x"090" => q <= x"00";
            when x"091" => q <= x"00";
            when x"092" => q <= x"00";
            when x"093" => q <= x"00";
            when x"094" => q <= x"00";
            when x"095" => q <= x"00";
            when x"096" => q <= x"00";
            when x"097" => q <= x"00";
            when x"098" => q <= x"00";
            when x"099" => q <= x"00";
            when x"09A" => q <= x"00";
            when x"09B" => q <= x"00";
            when x"09C" => q <= x"00";
            when x"09D" => q <= x"00";
            when x"09E" => q <= x"00";
            when x"09F" => q <= x"00";
            when x"0A0" => q <= x"00";
            when x"0A1" => q <= x"00";
            when x"0A2" => q <= x"00";
            when x"0A3" => q <= x"00";
            when x"0A4" => q <= x"00";
            when x"0A5" => q <= x"00";
            when x"0A6" => q <= x"00";
            when x"0A7" => q <= x"00";
            when x"0A8" => q <= x"00";
            when x"0A9" => q <= x"00";
            when x"0AA" => q <= x"00";
            when x"0AB" => q <= x"00";
            when x"0AC" => q <= x"00";
            when x"0AD" => q <= x"00";
            when x"0AE" => q <= x"00";
            when x"0AF" => q <= x"00";
            when x"0B0" => q <= x"00";
            when x"0B1" => q <= x"00";
            when x"0B2" => q <= x"00";
            when x"0B3" => q <= x"00";
            when x"0B4" => q <= x"00";
            when x"0B5" => q <= x"00";
            when x"0B6" => q <= x"00";
            when x"0B7" => q <= x"00";
            when x"0B8" => q <= x"00";
            when x"0B9" => q <= x"00";
            when x"0BA" => q <= x"00";
            when x"0BB" => q <= x"00";
            when x"0BC" => q <= x"00";
            when x"0BD" => q <= x"00";
            when x"0BE" => q <= x"00";
            when x"0BF" => q <= x"00";
            when x"0C0" => q <= x"00";
            when x"0C1" => q <= x"00";
            when x"0C2" => q <= x"00";
            when x"0C3" => q <= x"00";
            when x"0C4" => q <= x"00";
            when x"0C5" => q <= x"00";
            when x"0C6" => q <= x"00";
            when x"0C7" => q <= x"00";
            when x"0C8" => q <= x"00";
            when x"0C9" => q <= x"00";
            when x"0CA" => q <= x"00";
            when x"0CB" => q <= x"00";
            when x"0CC" => q <= x"00";
            when x"0CD" => q <= x"00";
            when x"0CE" => q <= x"00";
            when x"0CF" => q <= x"00";
            when x"0D0" => q <= x"00";
            when x"0D1" => q <= x"00";
            when x"0D2" => q <= x"00";
            when x"0D3" => q <= x"00";
            when x"0D4" => q <= x"00";
            when x"0D5" => q <= x"00";
            when x"0D6" => q <= x"00";
            when x"0D7" => q <= x"00";
            when x"0D8" => q <= x"00";
            when x"0D9" => q <= x"00";
            when x"0DA" => q <= x"00";
            when x"0DB" => q <= x"00";
            when x"0DC" => q <= x"00";
            when x"0DD" => q <= x"00";
            when x"0DE" => q <= x"00";
            when x"0DF" => q <= x"00";
            when x"0E0" => q <= x"00";
            when x"0E1" => q <= x"00";
            when x"0E2" => q <= x"00";
            when x"0E3" => q <= x"00";
            when x"0E4" => q <= x"00";
            when x"0E5" => q <= x"00";
            when x"0E6" => q <= x"00";
            when x"0E7" => q <= x"00";
            when x"0E8" => q <= x"00";
            when x"0E9" => q <= x"00";
            when x"0EA" => q <= x"00";
            when x"0EB" => q <= x"00";
            when x"0EC" => q <= x"00";
            when x"0ED" => q <= x"00";
            when x"0EE" => q <= x"00";
            when x"0EF" => q <= x"00";
            when x"0F0" => q <= x"00";
            when x"0F1" => q <= x"00";
            when x"0F2" => q <= x"00";
            when x"0F3" => q <= x"00";
            when x"0F4" => q <= x"00";
            when x"0F5" => q <= x"00";
            when x"0F6" => q <= x"00";
            when x"0F7" => q <= x"00";
            when x"0F8" => q <= x"00";
            when x"0F9" => q <= x"00";
            when x"0FA" => q <= x"00";
            when x"0FB" => q <= x"00";
            when x"0FC" => q <= x"00";
            when x"0FD" => q <= x"00";
            when x"0FE" => q <= x"00";
            when x"0FF" => q <= x"00";
            when x"100" => q <= x"00";
            when x"101" => q <= x"00";
            when x"102" => q <= x"00";
            when x"103" => q <= x"00";
            when x"104" => q <= x"00";
            when x"105" => q <= x"00";
            when x"106" => q <= x"00";
            when x"107" => q <= x"00";
            when x"108" => q <= x"00";
            when x"109" => q <= x"00";
            when x"10A" => q <= x"00";
            when x"10B" => q <= x"00";
            when x"10C" => q <= x"00";
            when x"10D" => q <= x"00";
            when x"10E" => q <= x"00";
            when x"10F" => q <= x"00";
            when x"110" => q <= x"00";
            when x"111" => q <= x"00";
            when x"112" => q <= x"00";
            when x"113" => q <= x"00";
            when x"114" => q <= x"00";
            when x"115" => q <= x"00";
            when x"116" => q <= x"00";
            when x"117" => q <= x"00";
            when x"118" => q <= x"00";
            when x"119" => q <= x"00";
            when x"11A" => q <= x"00";
            when x"11B" => q <= x"00";
            when x"11C" => q <= x"00";
            when x"11D" => q <= x"00";
            when x"11E" => q <= x"00";
            when x"11F" => q <= x"00";
            when x"120" => q <= x"00";
            when x"121" => q <= x"00";
            when x"122" => q <= x"00";
            when x"123" => q <= x"00";
            when x"124" => q <= x"00";
            when x"125" => q <= x"00";
            when x"126" => q <= x"00";
            when x"127" => q <= x"00";
            when x"128" => q <= x"00";
            when x"129" => q <= x"00";
            when x"12A" => q <= x"00";
            when x"12B" => q <= x"00";
            when x"12C" => q <= x"00";
            when x"12D" => q <= x"00";
            when x"12E" => q <= x"00";
            when x"12F" => q <= x"00";
            when x"130" => q <= x"00";
            when x"131" => q <= x"00";
            when x"132" => q <= x"00";
            when x"133" => q <= x"00";
            when x"134" => q <= x"00";
            when x"135" => q <= x"00";
            when x"136" => q <= x"00";
            when x"137" => q <= x"00";
            when x"138" => q <= x"00";
            when x"139" => q <= x"00";
            when x"13A" => q <= x"00";
            when x"13B" => q <= x"00";
            when x"13C" => q <= x"00";
            when x"13D" => q <= x"00";
            when x"13E" => q <= x"00";
            when x"13F" => q <= x"00";
            when x"140" => q <= x"00";
            when x"141" => q <= x"00";
            when x"142" => q <= x"00";
            when x"143" => q <= x"00";
            when x"144" => q <= x"00";
            when x"145" => q <= x"00";
            when x"146" => q <= x"00";
            when x"147" => q <= x"00";
            when x"148" => q <= x"00";
            when x"149" => q <= x"00";
            when x"14A" => q <= x"00";
            when x"14B" => q <= x"00";
            when x"14C" => q <= x"00";
            when x"14D" => q <= x"00";
            when x"14E" => q <= x"00";
            when x"14F" => q <= x"00";
            when x"150" => q <= x"00";
            when x"151" => q <= x"00";
            when x"152" => q <= x"00";
            when x"153" => q <= x"00";
            when x"154" => q <= x"00";
            when x"155" => q <= x"00";
            when x"156" => q <= x"00";
            when x"157" => q <= x"00";
            when x"158" => q <= x"00";
            when x"159" => q <= x"00";
            when x"15A" => q <= x"00";
            when x"15B" => q <= x"00";
            when x"15C" => q <= x"00";
            when x"15D" => q <= x"00";
            when x"15E" => q <= x"00";
            when x"15F" => q <= x"00";
            when x"160" => q <= x"00";
            when x"161" => q <= x"00";
            when x"162" => q <= x"00";
            when x"163" => q <= x"00";
            when x"164" => q <= x"00";
            when x"165" => q <= x"00";
            when x"166" => q <= x"00";
            when x"167" => q <= x"00";
            when x"168" => q <= x"00";
            when x"169" => q <= x"00";
            when x"16A" => q <= x"00";
            when x"16B" => q <= x"00";
            when x"16C" => q <= x"00";
            when x"16D" => q <= x"00";
            when x"16E" => q <= x"00";
            when x"16F" => q <= x"00";
            when x"170" => q <= x"00";
            when x"171" => q <= x"00";
            when x"172" => q <= x"00";
            when x"173" => q <= x"00";
            when x"174" => q <= x"00";
            when x"175" => q <= x"00";
            when x"176" => q <= x"00";
            when x"177" => q <= x"00";
            when x"178" => q <= x"00";
            when x"179" => q <= x"00";
            when x"17A" => q <= x"00";
            when x"17B" => q <= x"00";
            when x"17C" => q <= x"00";
            when x"17D" => q <= x"00";
            when x"17E" => q <= x"00";
            when x"17F" => q <= x"00";
            when x"180" => q <= x"00";
            when x"181" => q <= x"00";
            when x"182" => q <= x"00";
            when x"183" => q <= x"00";
            when x"184" => q <= x"00";
            when x"185" => q <= x"00";
            when x"186" => q <= x"00";
            when x"187" => q <= x"00";
            when x"188" => q <= x"00";
            when x"189" => q <= x"00";
            when x"18A" => q <= x"00";
            when x"18B" => q <= x"00";
            when x"18C" => q <= x"00";
            when x"18D" => q <= x"00";
            when x"18E" => q <= x"00";
            when x"18F" => q <= x"00";
            when x"190" => q <= x"00";
            when x"191" => q <= x"00";
            when x"192" => q <= x"00";
            when x"193" => q <= x"00";
            when x"194" => q <= x"00";
            when x"195" => q <= x"00";
            when x"196" => q <= x"00";
            when x"197" => q <= x"00";
            when x"198" => q <= x"00";
            when x"199" => q <= x"00";
            when x"19A" => q <= x"00";
            when x"19B" => q <= x"00";
            when x"19C" => q <= x"00";
            when x"19D" => q <= x"00";
            when x"19E" => q <= x"00";
            when x"19F" => q <= x"00";
            when x"1A0" => q <= x"00";
            when x"1A1" => q <= x"00";
            when x"1A2" => q <= x"00";
            when x"1A3" => q <= x"00";
            when x"1A4" => q <= x"00";
            when x"1A5" => q <= x"00";
            when x"1A6" => q <= x"00";
            when x"1A7" => q <= x"00";
            when x"1A8" => q <= x"00";
            when x"1A9" => q <= x"00";
            when x"1AA" => q <= x"00";
            when x"1AB" => q <= x"00";
            when x"1AC" => q <= x"00";
            when x"1AD" => q <= x"00";
            when x"1AE" => q <= x"00";
            when x"1AF" => q <= x"00";
            when x"1B0" => q <= x"00";
            when x"1B1" => q <= x"00";
            when x"1B2" => q <= x"00";
            when x"1B3" => q <= x"00";
            when x"1B4" => q <= x"00";
            when x"1B5" => q <= x"00";
            when x"1B6" => q <= x"00";
            when x"1B7" => q <= x"00";
            when x"1B8" => q <= x"00";
            when x"1B9" => q <= x"00";
            when x"1BA" => q <= x"00";
            when x"1BB" => q <= x"00";
            when x"1BC" => q <= x"00";
            when x"1BD" => q <= x"00";
            when x"1BE" => q <= x"00";
            when x"1BF" => q <= x"00";
            when x"1C0" => q <= x"00";
            when x"1C1" => q <= x"00";
            when x"1C2" => q <= x"00";
            when x"1C3" => q <= x"00";
            when x"1C4" => q <= x"00";
            when x"1C5" => q <= x"00";
            when x"1C6" => q <= x"00";
            when x"1C7" => q <= x"00";
            when x"1C8" => q <= x"00";
            when x"1C9" => q <= x"00";
            when x"1CA" => q <= x"00";
            when x"1CB" => q <= x"00";
            when x"1CC" => q <= x"00";
            when x"1CD" => q <= x"00";
            when x"1CE" => q <= x"00";
            when x"1CF" => q <= x"00";
            when x"1D0" => q <= x"00";
            when x"1D1" => q <= x"00";
            when x"1D2" => q <= x"00";
            when x"1D3" => q <= x"00";
            when x"1D4" => q <= x"00";
            when x"1D5" => q <= x"00";
            when x"1D6" => q <= x"00";
            when x"1D7" => q <= x"00";
            when x"1D8" => q <= x"00";
            when x"1D9" => q <= x"00";
            when x"1DA" => q <= x"00";
            when x"1DB" => q <= x"00";
            when x"1DC" => q <= x"00";
            when x"1DD" => q <= x"00";
            when x"1DE" => q <= x"00";
            when x"1DF" => q <= x"00";
            when x"1E0" => q <= x"00";
            when x"1E1" => q <= x"00";
            when x"1E2" => q <= x"00";
            when x"1E3" => q <= x"00";
            when x"1E4" => q <= x"00";
            when x"1E5" => q <= x"00";
            when x"1E6" => q <= x"00";
            when x"1E7" => q <= x"00";
            when x"1E8" => q <= x"00";
            when x"1E9" => q <= x"00";
            when x"1EA" => q <= x"00";
            when x"1EB" => q <= x"00";
            when x"1EC" => q <= x"00";
            when x"1ED" => q <= x"00";
            when x"1EE" => q <= x"00";
            when x"1EF" => q <= x"00";
            when x"1F0" => q <= x"00";
            when x"1F1" => q <= x"00";
            when x"1F2" => q <= x"00";
            when x"1F3" => q <= x"00";
            when x"1F4" => q <= x"00";
            when x"1F5" => q <= x"00";
            when x"1F6" => q <= x"00";
            when x"1F7" => q <= x"00";
            when x"1F8" => q <= x"00";
            when x"1F9" => q <= x"00";
            when x"1FA" => q <= x"00";
            when x"1FB" => q <= x"00";
            when x"1FC" => q <= x"00";
            when x"1FD" => q <= x"00";
            when x"1FE" => q <= x"00";
            when x"1FF" => q <= x"00";
            when x"200" => q <= x"00";
            when x"201" => q <= x"00";
            when x"202" => q <= x"00";
            when x"203" => q <= x"00";
            when x"204" => q <= x"00";
            when x"205" => q <= x"00";
            when x"206" => q <= x"00";
            when x"207" => q <= x"00";
            when x"208" => q <= x"00";
            when x"209" => q <= x"00";
            when x"20A" => q <= x"00";
            when x"20B" => q <= x"00";
            when x"20C" => q <= x"00";
            when x"20D" => q <= x"00";
            when x"20E" => q <= x"00";
            when x"20F" => q <= x"00";
            when x"210" => q <= x"00";
            when x"211" => q <= x"04";
            when x"212" => q <= x"04";
            when x"213" => q <= x"04";
            when x"214" => q <= x"04";
            when x"215" => q <= x"04";
            when x"216" => q <= x"00";
            when x"217" => q <= x"04";
            when x"218" => q <= x"00";
            when x"219" => q <= x"00";
            when x"21A" => q <= x"00";
            when x"21B" => q <= x"00";
            when x"21C" => q <= x"00";
            when x"21D" => q <= x"00";
            when x"21E" => q <= x"00";
            when x"21F" => q <= x"00";
            when x"220" => q <= x"00";
            when x"221" => q <= x"0A";
            when x"222" => q <= x"0A";
            when x"223" => q <= x"0A";
            when x"224" => q <= x"00";
            when x"225" => q <= x"00";
            when x"226" => q <= x"00";
            when x"227" => q <= x"00";
            when x"228" => q <= x"00";
            when x"229" => q <= x"00";
            when x"22A" => q <= x"00";
            when x"22B" => q <= x"00";
            when x"22C" => q <= x"00";
            when x"22D" => q <= x"00";
            when x"22E" => q <= x"00";
            when x"22F" => q <= x"00";
            when x"230" => q <= x"00";
            when x"231" => q <= x"06";
            when x"232" => q <= x"09";
            when x"233" => q <= x"08";
            when x"234" => q <= x"1C";
            when x"235" => q <= x"08";
            when x"236" => q <= x"08";
            when x"237" => q <= x"1F";
            when x"238" => q <= x"00";
            when x"239" => q <= x"00";
            when x"23A" => q <= x"00";
            when x"23B" => q <= x"00";
            when x"23C" => q <= x"00";
            when x"23D" => q <= x"00";
            when x"23E" => q <= x"00";
            when x"23F" => q <= x"00";
            when x"240" => q <= x"00";
            when x"241" => q <= x"0E";
            when x"242" => q <= x"15";
            when x"243" => q <= x"14";
            when x"244" => q <= x"0E";
            when x"245" => q <= x"05";
            when x"246" => q <= x"15";
            when x"247" => q <= x"0E";
            when x"248" => q <= x"00";
            when x"249" => q <= x"00";
            when x"24A" => q <= x"00";
            when x"24B" => q <= x"00";
            when x"24C" => q <= x"00";
            when x"24D" => q <= x"00";
            when x"24E" => q <= x"00";
            when x"24F" => q <= x"00";
            when x"250" => q <= x"00";
            when x"251" => q <= x"18";
            when x"252" => q <= x"19";
            when x"253" => q <= x"02";
            when x"254" => q <= x"04";
            when x"255" => q <= x"08";
            when x"256" => q <= x"13";
            when x"257" => q <= x"03";
            when x"258" => q <= x"00";
            when x"259" => q <= x"00";
            when x"25A" => q <= x"00";
            when x"25B" => q <= x"00";
            when x"25C" => q <= x"00";
            when x"25D" => q <= x"00";
            when x"25E" => q <= x"00";
            when x"25F" => q <= x"00";
            when x"260" => q <= x"00";
            when x"261" => q <= x"08";
            when x"262" => q <= x"14";
            when x"263" => q <= x"14";
            when x"264" => q <= x"08";
            when x"265" => q <= x"15";
            when x"266" => q <= x"12";
            when x"267" => q <= x"0D";
            when x"268" => q <= x"00";
            when x"269" => q <= x"00";
            when x"26A" => q <= x"00";
            when x"26B" => q <= x"00";
            when x"26C" => q <= x"00";
            when x"26D" => q <= x"00";
            when x"26E" => q <= x"00";
            when x"26F" => q <= x"00";
            when x"270" => q <= x"00";
            when x"271" => q <= x"04";
            when x"272" => q <= x"04";
            when x"273" => q <= x"04";
            when x"274" => q <= x"00";
            when x"275" => q <= x"00";
            when x"276" => q <= x"00";
            when x"277" => q <= x"00";
            when x"278" => q <= x"00";
            when x"279" => q <= x"00";
            when x"27A" => q <= x"00";
            when x"27B" => q <= x"00";
            when x"27C" => q <= x"00";
            when x"27D" => q <= x"00";
            when x"27E" => q <= x"00";
            when x"27F" => q <= x"00";
            when x"280" => q <= x"00";
            when x"281" => q <= x"02";
            when x"282" => q <= x"04";
            when x"283" => q <= x"08";
            when x"284" => q <= x"08";
            when x"285" => q <= x"08";
            when x"286" => q <= x"04";
            when x"287" => q <= x"02";
            when x"288" => q <= x"00";
            when x"289" => q <= x"00";
            when x"28A" => q <= x"00";
            when x"28B" => q <= x"00";
            when x"28C" => q <= x"00";
            when x"28D" => q <= x"00";
            when x"28E" => q <= x"00";
            when x"28F" => q <= x"00";
            when x"290" => q <= x"00";
            when x"291" => q <= x"08";
            when x"292" => q <= x"04";
            when x"293" => q <= x"02";
            when x"294" => q <= x"02";
            when x"295" => q <= x"02";
            when x"296" => q <= x"04";
            when x"297" => q <= x"08";
            when x"298" => q <= x"00";
            when x"299" => q <= x"00";
            when x"29A" => q <= x"00";
            when x"29B" => q <= x"00";
            when x"29C" => q <= x"00";
            when x"29D" => q <= x"00";
            when x"29E" => q <= x"00";
            when x"29F" => q <= x"00";
            when x"2A0" => q <= x"00";
            when x"2A1" => q <= x"04";
            when x"2A2" => q <= x"15";
            when x"2A3" => q <= x"0E";
            when x"2A4" => q <= x"04";
            when x"2A5" => q <= x"0E";
            when x"2A6" => q <= x"15";
            when x"2A7" => q <= x"04";
            when x"2A8" => q <= x"00";
            when x"2A9" => q <= x"00";
            when x"2AA" => q <= x"00";
            when x"2AB" => q <= x"00";
            when x"2AC" => q <= x"00";
            when x"2AD" => q <= x"00";
            when x"2AE" => q <= x"00";
            when x"2AF" => q <= x"00";
            when x"2B0" => q <= x"00";
            when x"2B1" => q <= x"00";
            when x"2B2" => q <= x"04";
            when x"2B3" => q <= x"04";
            when x"2B4" => q <= x"1F";
            when x"2B5" => q <= x"04";
            when x"2B6" => q <= x"04";
            when x"2B7" => q <= x"00";
            when x"2B8" => q <= x"00";
            when x"2B9" => q <= x"00";
            when x"2BA" => q <= x"00";
            when x"2BB" => q <= x"00";
            when x"2BC" => q <= x"00";
            when x"2BD" => q <= x"00";
            when x"2BE" => q <= x"00";
            when x"2BF" => q <= x"00";
            when x"2C0" => q <= x"00";
            when x"2C1" => q <= x"00";
            when x"2C2" => q <= x"00";
            when x"2C3" => q <= x"00";
            when x"2C4" => q <= x"00";
            when x"2C5" => q <= x"00";
            when x"2C6" => q <= x"04";
            when x"2C7" => q <= x"04";
            when x"2C8" => q <= x"08";
            when x"2C9" => q <= x"00";
            when x"2CA" => q <= x"00";
            when x"2CB" => q <= x"00";
            when x"2CC" => q <= x"00";
            when x"2CD" => q <= x"00";
            when x"2CE" => q <= x"00";
            when x"2CF" => q <= x"00";
            when x"2D0" => q <= x"00";
            when x"2D1" => q <= x"00";
            when x"2D2" => q <= x"00";
            when x"2D3" => q <= x"00";
            when x"2D4" => q <= x"0E";
            when x"2D5" => q <= x"00";
            when x"2D6" => q <= x"00";
            when x"2D7" => q <= x"00";
            when x"2D8" => q <= x"00";
            when x"2D9" => q <= x"00";
            when x"2DA" => q <= x"00";
            when x"2DB" => q <= x"00";
            when x"2DC" => q <= x"00";
            when x"2DD" => q <= x"00";
            when x"2DE" => q <= x"00";
            when x"2DF" => q <= x"00";
            when x"2E0" => q <= x"00";
            when x"2E1" => q <= x"00";
            when x"2E2" => q <= x"00";
            when x"2E3" => q <= x"00";
            when x"2E4" => q <= x"00";
            when x"2E5" => q <= x"00";
            when x"2E6" => q <= x"00";
            when x"2E7" => q <= x"04";
            when x"2E8" => q <= x"00";
            when x"2E9" => q <= x"00";
            when x"2EA" => q <= x"00";
            when x"2EB" => q <= x"00";
            when x"2EC" => q <= x"00";
            when x"2ED" => q <= x"00";
            when x"2EE" => q <= x"00";
            when x"2EF" => q <= x"00";
            when x"2F0" => q <= x"00";
            when x"2F1" => q <= x"00";
            when x"2F2" => q <= x"01";
            when x"2F3" => q <= x"02";
            when x"2F4" => q <= x"04";
            when x"2F5" => q <= x"08";
            when x"2F6" => q <= x"10";
            when x"2F7" => q <= x"00";
            when x"2F8" => q <= x"00";
            when x"2F9" => q <= x"00";
            when x"2FA" => q <= x"00";
            when x"2FB" => q <= x"00";
            when x"2FC" => q <= x"00";
            when x"2FD" => q <= x"00";
            when x"2FE" => q <= x"00";
            when x"2FF" => q <= x"00";
            when x"300" => q <= x"00";
            when x"301" => q <= x"04";
            when x"302" => q <= x"0A";
            when x"303" => q <= x"11";
            when x"304" => q <= x"11";
            when x"305" => q <= x"11";
            when x"306" => q <= x"0A";
            when x"307" => q <= x"04";
            when x"308" => q <= x"00";
            when x"309" => q <= x"00";
            when x"30A" => q <= x"00";
            when x"30B" => q <= x"00";
            when x"30C" => q <= x"00";
            when x"30D" => q <= x"00";
            when x"30E" => q <= x"00";
            when x"30F" => q <= x"00";
            when x"310" => q <= x"00";
            when x"311" => q <= x"04";
            when x"312" => q <= x"0C";
            when x"313" => q <= x"04";
            when x"314" => q <= x"04";
            when x"315" => q <= x"04";
            when x"316" => q <= x"04";
            when x"317" => q <= x"0E";
            when x"318" => q <= x"00";
            when x"319" => q <= x"00";
            when x"31A" => q <= x"00";
            when x"31B" => q <= x"00";
            when x"31C" => q <= x"00";
            when x"31D" => q <= x"00";
            when x"31E" => q <= x"00";
            when x"31F" => q <= x"00";
            when x"320" => q <= x"00";
            when x"321" => q <= x"0E";
            when x"322" => q <= x"11";
            when x"323" => q <= x"01";
            when x"324" => q <= x"06";
            when x"325" => q <= x"08";
            when x"326" => q <= x"10";
            when x"327" => q <= x"1F";
            when x"328" => q <= x"00";
            when x"329" => q <= x"00";
            when x"32A" => q <= x"00";
            when x"32B" => q <= x"00";
            when x"32C" => q <= x"00";
            when x"32D" => q <= x"00";
            when x"32E" => q <= x"00";
            when x"32F" => q <= x"00";
            when x"330" => q <= x"00";
            when x"331" => q <= x"1F";
            when x"332" => q <= x"01";
            when x"333" => q <= x"02";
            when x"334" => q <= x"06";
            when x"335" => q <= x"01";
            when x"336" => q <= x"11";
            when x"337" => q <= x"0E";
            when x"338" => q <= x"00";
            when x"339" => q <= x"00";
            when x"33A" => q <= x"00";
            when x"33B" => q <= x"00";
            when x"33C" => q <= x"00";
            when x"33D" => q <= x"00";
            when x"33E" => q <= x"00";
            when x"33F" => q <= x"00";
            when x"340" => q <= x"00";
            when x"341" => q <= x"02";
            when x"342" => q <= x"06";
            when x"343" => q <= x"0A";
            when x"344" => q <= x"12";
            when x"345" => q <= x"1F";
            when x"346" => q <= x"02";
            when x"347" => q <= x"02";
            when x"348" => q <= x"00";
            when x"349" => q <= x"00";
            when x"34A" => q <= x"00";
            when x"34B" => q <= x"00";
            when x"34C" => q <= x"00";
            when x"34D" => q <= x"00";
            when x"34E" => q <= x"00";
            when x"34F" => q <= x"00";
            when x"350" => q <= x"00";
            when x"351" => q <= x"1F";
            when x"352" => q <= x"10";
            when x"353" => q <= x"1E";
            when x"354" => q <= x"01";
            when x"355" => q <= x"01";
            when x"356" => q <= x"11";
            when x"357" => q <= x"0E";
            when x"358" => q <= x"00";
            when x"359" => q <= x"00";
            when x"35A" => q <= x"00";
            when x"35B" => q <= x"00";
            when x"35C" => q <= x"00";
            when x"35D" => q <= x"00";
            when x"35E" => q <= x"00";
            when x"35F" => q <= x"00";
            when x"360" => q <= x"00";
            when x"361" => q <= x"06";
            when x"362" => q <= x"08";
            when x"363" => q <= x"10";
            when x"364" => q <= x"1E";
            when x"365" => q <= x"11";
            when x"366" => q <= x"11";
            when x"367" => q <= x"0E";
            when x"368" => q <= x"00";
            when x"369" => q <= x"00";
            when x"36A" => q <= x"00";
            when x"36B" => q <= x"00";
            when x"36C" => q <= x"00";
            when x"36D" => q <= x"00";
            when x"36E" => q <= x"00";
            when x"36F" => q <= x"00";
            when x"370" => q <= x"00";
            when x"371" => q <= x"1F";
            when x"372" => q <= x"01";
            when x"373" => q <= x"02";
            when x"374" => q <= x"04";
            when x"375" => q <= x"08";
            when x"376" => q <= x"08";
            when x"377" => q <= x"08";
            when x"378" => q <= x"00";
            when x"379" => q <= x"00";
            when x"37A" => q <= x"00";
            when x"37B" => q <= x"00";
            when x"37C" => q <= x"00";
            when x"37D" => q <= x"00";
            when x"37E" => q <= x"00";
            when x"37F" => q <= x"00";
            when x"380" => q <= x"00";
            when x"381" => q <= x"0E";
            when x"382" => q <= x"11";
            when x"383" => q <= x"11";
            when x"384" => q <= x"0E";
            when x"385" => q <= x"11";
            when x"386" => q <= x"11";
            when x"387" => q <= x"0E";
            when x"388" => q <= x"00";
            when x"389" => q <= x"00";
            when x"38A" => q <= x"00";
            when x"38B" => q <= x"00";
            when x"38C" => q <= x"00";
            when x"38D" => q <= x"00";
            when x"38E" => q <= x"00";
            when x"38F" => q <= x"00";
            when x"390" => q <= x"00";
            when x"391" => q <= x"0E";
            when x"392" => q <= x"11";
            when x"393" => q <= x"11";
            when x"394" => q <= x"0F";
            when x"395" => q <= x"01";
            when x"396" => q <= x"02";
            when x"397" => q <= x"0C";
            when x"398" => q <= x"00";
            when x"399" => q <= x"00";
            when x"39A" => q <= x"00";
            when x"39B" => q <= x"00";
            when x"39C" => q <= x"00";
            when x"39D" => q <= x"00";
            when x"39E" => q <= x"00";
            when x"39F" => q <= x"00";
            when x"3A0" => q <= x"00";
            when x"3A1" => q <= x"00";
            when x"3A2" => q <= x"00";
            when x"3A3" => q <= x"04";
            when x"3A4" => q <= x"00";
            when x"3A5" => q <= x"00";
            when x"3A6" => q <= x"00";
            when x"3A7" => q <= x"04";
            when x"3A8" => q <= x"00";
            when x"3A9" => q <= x"00";
            when x"3AA" => q <= x"00";
            when x"3AB" => q <= x"00";
            when x"3AC" => q <= x"00";
            when x"3AD" => q <= x"00";
            when x"3AE" => q <= x"00";
            when x"3AF" => q <= x"00";
            when x"3B0" => q <= x"00";
            when x"3B1" => q <= x"00";
            when x"3B2" => q <= x"00";
            when x"3B3" => q <= x"04";
            when x"3B4" => q <= x"00";
            when x"3B5" => q <= x"00";
            when x"3B6" => q <= x"04";
            when x"3B7" => q <= x"04";
            when x"3B8" => q <= x"08";
            when x"3B9" => q <= x"00";
            when x"3BA" => q <= x"00";
            when x"3BB" => q <= x"00";
            when x"3BC" => q <= x"00";
            when x"3BD" => q <= x"00";
            when x"3BE" => q <= x"00";
            when x"3BF" => q <= x"00";
            when x"3C0" => q <= x"00";
            when x"3C1" => q <= x"02";
            when x"3C2" => q <= x"04";
            when x"3C3" => q <= x"08";
            when x"3C4" => q <= x"10";
            when x"3C5" => q <= x"08";
            when x"3C6" => q <= x"04";
            when x"3C7" => q <= x"02";
            when x"3C8" => q <= x"00";
            when x"3C9" => q <= x"00";
            when x"3CA" => q <= x"00";
            when x"3CB" => q <= x"00";
            when x"3CC" => q <= x"00";
            when x"3CD" => q <= x"00";
            when x"3CE" => q <= x"00";
            when x"3CF" => q <= x"00";
            when x"3D0" => q <= x"00";
            when x"3D1" => q <= x"00";
            when x"3D2" => q <= x"00";
            when x"3D3" => q <= x"1F";
            when x"3D4" => q <= x"00";
            when x"3D5" => q <= x"1F";
            when x"3D6" => q <= x"00";
            when x"3D7" => q <= x"00";
            when x"3D8" => q <= x"00";
            when x"3D9" => q <= x"00";
            when x"3DA" => q <= x"00";
            when x"3DB" => q <= x"00";
            when x"3DC" => q <= x"00";
            when x"3DD" => q <= x"00";
            when x"3DE" => q <= x"00";
            when x"3DF" => q <= x"00";
            when x"3E0" => q <= x"00";
            when x"3E1" => q <= x"08";
            when x"3E2" => q <= x"04";
            when x"3E3" => q <= x"02";
            when x"3E4" => q <= x"01";
            when x"3E5" => q <= x"02";
            when x"3E6" => q <= x"04";
            when x"3E7" => q <= x"08";
            when x"3E8" => q <= x"00";
            when x"3E9" => q <= x"00";
            when x"3EA" => q <= x"00";
            when x"3EB" => q <= x"00";
            when x"3EC" => q <= x"00";
            when x"3ED" => q <= x"00";
            when x"3EE" => q <= x"00";
            when x"3EF" => q <= x"00";
            when x"3F0" => q <= x"00";
            when x"3F1" => q <= x"0E";
            when x"3F2" => q <= x"11";
            when x"3F3" => q <= x"02";
            when x"3F4" => q <= x"04";
            when x"3F5" => q <= x"04";
            when x"3F6" => q <= x"00";
            when x"3F7" => q <= x"04";
            when x"3F8" => q <= x"00";
            when x"3F9" => q <= x"00";
            when x"3FA" => q <= x"00";
            when x"3FB" => q <= x"00";
            when x"3FC" => q <= x"00";
            when x"3FD" => q <= x"00";
            when x"3FE" => q <= x"00";
            when x"3FF" => q <= x"00";
            when x"400" => q <= x"00";
            when x"401" => q <= x"0E";
            when x"402" => q <= x"11";
            when x"403" => q <= x"17";
            when x"404" => q <= x"15";
            when x"405" => q <= x"17";
            when x"406" => q <= x"10";
            when x"407" => q <= x"0E";
            when x"408" => q <= x"00";
            when x"409" => q <= x"00";
            when x"40A" => q <= x"00";
            when x"40B" => q <= x"00";
            when x"40C" => q <= x"00";
            when x"40D" => q <= x"00";
            when x"40E" => q <= x"00";
            when x"40F" => q <= x"00";
            when x"410" => q <= x"00";
            when x"411" => q <= x"04";
            when x"412" => q <= x"0A";
            when x"413" => q <= x"11";
            when x"414" => q <= x"11";
            when x"415" => q <= x"1F";
            when x"416" => q <= x"11";
            when x"417" => q <= x"11";
            when x"418" => q <= x"00";
            when x"419" => q <= x"00";
            when x"41A" => q <= x"00";
            when x"41B" => q <= x"00";
            when x"41C" => q <= x"00";
            when x"41D" => q <= x"00";
            when x"41E" => q <= x"00";
            when x"41F" => q <= x"00";
            when x"420" => q <= x"00";
            when x"421" => q <= x"1E";
            when x"422" => q <= x"11";
            when x"423" => q <= x"11";
            when x"424" => q <= x"1E";
            when x"425" => q <= x"11";
            when x"426" => q <= x"11";
            when x"427" => q <= x"1E";
            when x"428" => q <= x"00";
            when x"429" => q <= x"00";
            when x"42A" => q <= x"00";
            when x"42B" => q <= x"00";
            when x"42C" => q <= x"00";
            when x"42D" => q <= x"00";
            when x"42E" => q <= x"00";
            when x"42F" => q <= x"00";
            when x"430" => q <= x"00";
            when x"431" => q <= x"0E";
            when x"432" => q <= x"11";
            when x"433" => q <= x"10";
            when x"434" => q <= x"10";
            when x"435" => q <= x"10";
            when x"436" => q <= x"11";
            when x"437" => q <= x"0E";
            when x"438" => q <= x"00";
            when x"439" => q <= x"00";
            when x"43A" => q <= x"00";
            when x"43B" => q <= x"00";
            when x"43C" => q <= x"00";
            when x"43D" => q <= x"00";
            when x"43E" => q <= x"00";
            when x"43F" => q <= x"00";
            when x"440" => q <= x"00";
            when x"441" => q <= x"1E";
            when x"442" => q <= x"11";
            when x"443" => q <= x"11";
            when x"444" => q <= x"11";
            when x"445" => q <= x"11";
            when x"446" => q <= x"11";
            when x"447" => q <= x"1E";
            when x"448" => q <= x"00";
            when x"449" => q <= x"00";
            when x"44A" => q <= x"00";
            when x"44B" => q <= x"00";
            when x"44C" => q <= x"00";
            when x"44D" => q <= x"00";
            when x"44E" => q <= x"00";
            when x"44F" => q <= x"00";
            when x"450" => q <= x"00";
            when x"451" => q <= x"1F";
            when x"452" => q <= x"10";
            when x"453" => q <= x"10";
            when x"454" => q <= x"1E";
            when x"455" => q <= x"10";
            when x"456" => q <= x"10";
            when x"457" => q <= x"1F";
            when x"458" => q <= x"00";
            when x"459" => q <= x"00";
            when x"45A" => q <= x"00";
            when x"45B" => q <= x"00";
            when x"45C" => q <= x"00";
            when x"45D" => q <= x"00";
            when x"45E" => q <= x"00";
            when x"45F" => q <= x"00";
            when x"460" => q <= x"00";
            when x"461" => q <= x"1F";
            when x"462" => q <= x"10";
            when x"463" => q <= x"10";
            when x"464" => q <= x"1E";
            when x"465" => q <= x"10";
            when x"466" => q <= x"10";
            when x"467" => q <= x"10";
            when x"468" => q <= x"00";
            when x"469" => q <= x"00";
            when x"46A" => q <= x"00";
            when x"46B" => q <= x"00";
            when x"46C" => q <= x"00";
            when x"46D" => q <= x"00";
            when x"46E" => q <= x"00";
            when x"46F" => q <= x"00";
            when x"470" => q <= x"00";
            when x"471" => q <= x"0E";
            when x"472" => q <= x"11";
            when x"473" => q <= x"10";
            when x"474" => q <= x"10";
            when x"475" => q <= x"13";
            when x"476" => q <= x"11";
            when x"477" => q <= x"0F";
            when x"478" => q <= x"00";
            when x"479" => q <= x"00";
            when x"47A" => q <= x"00";
            when x"47B" => q <= x"00";
            when x"47C" => q <= x"00";
            when x"47D" => q <= x"00";
            when x"47E" => q <= x"00";
            when x"47F" => q <= x"00";
            when x"480" => q <= x"00";
            when x"481" => q <= x"11";
            when x"482" => q <= x"11";
            when x"483" => q <= x"11";
            when x"484" => q <= x"1F";
            when x"485" => q <= x"11";
            when x"486" => q <= x"11";
            when x"487" => q <= x"11";
            when x"488" => q <= x"00";
            when x"489" => q <= x"00";
            when x"48A" => q <= x"00";
            when x"48B" => q <= x"00";
            when x"48C" => q <= x"00";
            when x"48D" => q <= x"00";
            when x"48E" => q <= x"00";
            when x"48F" => q <= x"00";
            when x"490" => q <= x"00";
            when x"491" => q <= x"0E";
            when x"492" => q <= x"04";
            when x"493" => q <= x"04";
            when x"494" => q <= x"04";
            when x"495" => q <= x"04";
            when x"496" => q <= x"04";
            when x"497" => q <= x"0E";
            when x"498" => q <= x"00";
            when x"499" => q <= x"00";
            when x"49A" => q <= x"00";
            when x"49B" => q <= x"00";
            when x"49C" => q <= x"00";
            when x"49D" => q <= x"00";
            when x"49E" => q <= x"00";
            when x"49F" => q <= x"00";
            when x"4A0" => q <= x"00";
            when x"4A1" => q <= x"01";
            when x"4A2" => q <= x"01";
            when x"4A3" => q <= x"01";
            when x"4A4" => q <= x"01";
            when x"4A5" => q <= x"01";
            when x"4A6" => q <= x"11";
            when x"4A7" => q <= x"0E";
            when x"4A8" => q <= x"00";
            when x"4A9" => q <= x"00";
            when x"4AA" => q <= x"00";
            when x"4AB" => q <= x"00";
            when x"4AC" => q <= x"00";
            when x"4AD" => q <= x"00";
            when x"4AE" => q <= x"00";
            when x"4AF" => q <= x"00";
            when x"4B0" => q <= x"00";
            when x"4B1" => q <= x"11";
            when x"4B2" => q <= x"12";
            when x"4B3" => q <= x"14";
            when x"4B4" => q <= x"18";
            when x"4B5" => q <= x"14";
            when x"4B6" => q <= x"12";
            when x"4B7" => q <= x"11";
            when x"4B8" => q <= x"00";
            when x"4B9" => q <= x"00";
            when x"4BA" => q <= x"00";
            when x"4BB" => q <= x"00";
            when x"4BC" => q <= x"00";
            when x"4BD" => q <= x"00";
            when x"4BE" => q <= x"00";
            when x"4BF" => q <= x"00";
            when x"4C0" => q <= x"00";
            when x"4C1" => q <= x"10";
            when x"4C2" => q <= x"10";
            when x"4C3" => q <= x"10";
            when x"4C4" => q <= x"10";
            when x"4C5" => q <= x"10";
            when x"4C6" => q <= x"10";
            when x"4C7" => q <= x"1F";
            when x"4C8" => q <= x"00";
            when x"4C9" => q <= x"00";
            when x"4CA" => q <= x"00";
            when x"4CB" => q <= x"00";
            when x"4CC" => q <= x"00";
            when x"4CD" => q <= x"00";
            when x"4CE" => q <= x"00";
            when x"4CF" => q <= x"00";
            when x"4D0" => q <= x"00";
            when x"4D1" => q <= x"11";
            when x"4D2" => q <= x"1B";
            when x"4D3" => q <= x"15";
            when x"4D4" => q <= x"15";
            when x"4D5" => q <= x"11";
            when x"4D6" => q <= x"11";
            when x"4D7" => q <= x"11";
            when x"4D8" => q <= x"00";
            when x"4D9" => q <= x"00";
            when x"4DA" => q <= x"00";
            when x"4DB" => q <= x"00";
            when x"4DC" => q <= x"00";
            when x"4DD" => q <= x"00";
            when x"4DE" => q <= x"00";
            when x"4DF" => q <= x"00";
            when x"4E0" => q <= x"00";
            when x"4E1" => q <= x"11";
            when x"4E2" => q <= x"11";
            when x"4E3" => q <= x"19";
            when x"4E4" => q <= x"15";
            when x"4E5" => q <= x"13";
            when x"4E6" => q <= x"11";
            when x"4E7" => q <= x"11";
            when x"4E8" => q <= x"00";
            when x"4E9" => q <= x"00";
            when x"4EA" => q <= x"00";
            when x"4EB" => q <= x"00";
            when x"4EC" => q <= x"00";
            when x"4ED" => q <= x"00";
            when x"4EE" => q <= x"00";
            when x"4EF" => q <= x"00";
            when x"4F0" => q <= x"00";
            when x"4F1" => q <= x"0E";
            when x"4F2" => q <= x"11";
            when x"4F3" => q <= x"11";
            when x"4F4" => q <= x"11";
            when x"4F5" => q <= x"11";
            when x"4F6" => q <= x"11";
            when x"4F7" => q <= x"0E";
            when x"4F8" => q <= x"00";
            when x"4F9" => q <= x"00";
            when x"4FA" => q <= x"00";
            when x"4FB" => q <= x"00";
            when x"4FC" => q <= x"00";
            when x"4FD" => q <= x"00";
            when x"4FE" => q <= x"00";
            when x"4FF" => q <= x"00";
            when x"500" => q <= x"00";
            when x"501" => q <= x"1E";
            when x"502" => q <= x"11";
            when x"503" => q <= x"11";
            when x"504" => q <= x"1E";
            when x"505" => q <= x"10";
            when x"506" => q <= x"10";
            when x"507" => q <= x"10";
            when x"508" => q <= x"00";
            when x"509" => q <= x"00";
            when x"50A" => q <= x"00";
            when x"50B" => q <= x"00";
            when x"50C" => q <= x"00";
            when x"50D" => q <= x"00";
            when x"50E" => q <= x"00";
            when x"50F" => q <= x"00";
            when x"510" => q <= x"00";
            when x"511" => q <= x"0E";
            when x"512" => q <= x"11";
            when x"513" => q <= x"11";
            when x"514" => q <= x"11";
            when x"515" => q <= x"15";
            when x"516" => q <= x"12";
            when x"517" => q <= x"0D";
            when x"518" => q <= x"00";
            when x"519" => q <= x"00";
            when x"51A" => q <= x"00";
            when x"51B" => q <= x"00";
            when x"51C" => q <= x"00";
            when x"51D" => q <= x"00";
            when x"51E" => q <= x"00";
            when x"51F" => q <= x"00";
            when x"520" => q <= x"00";
            when x"521" => q <= x"1E";
            when x"522" => q <= x"11";
            when x"523" => q <= x"11";
            when x"524" => q <= x"1E";
            when x"525" => q <= x"14";
            when x"526" => q <= x"12";
            when x"527" => q <= x"11";
            when x"528" => q <= x"00";
            when x"529" => q <= x"00";
            when x"52A" => q <= x"00";
            when x"52B" => q <= x"00";
            when x"52C" => q <= x"00";
            when x"52D" => q <= x"00";
            when x"52E" => q <= x"00";
            when x"52F" => q <= x"00";
            when x"530" => q <= x"00";
            when x"531" => q <= x"0E";
            when x"532" => q <= x"11";
            when x"533" => q <= x"10";
            when x"534" => q <= x"0E";
            when x"535" => q <= x"01";
            when x"536" => q <= x"11";
            when x"537" => q <= x"0E";
            when x"538" => q <= x"00";
            when x"539" => q <= x"00";
            when x"53A" => q <= x"00";
            when x"53B" => q <= x"00";
            when x"53C" => q <= x"00";
            when x"53D" => q <= x"00";
            when x"53E" => q <= x"00";
            when x"53F" => q <= x"00";
            when x"540" => q <= x"00";
            when x"541" => q <= x"1F";
            when x"542" => q <= x"04";
            when x"543" => q <= x"04";
            when x"544" => q <= x"04";
            when x"545" => q <= x"04";
            when x"546" => q <= x"04";
            when x"547" => q <= x"04";
            when x"548" => q <= x"00";
            when x"549" => q <= x"00";
            when x"54A" => q <= x"00";
            when x"54B" => q <= x"00";
            when x"54C" => q <= x"00";
            when x"54D" => q <= x"00";
            when x"54E" => q <= x"00";
            when x"54F" => q <= x"00";
            when x"550" => q <= x"00";
            when x"551" => q <= x"11";
            when x"552" => q <= x"11";
            when x"553" => q <= x"11";
            when x"554" => q <= x"11";
            when x"555" => q <= x"11";
            when x"556" => q <= x"11";
            when x"557" => q <= x"0E";
            when x"558" => q <= x"00";
            when x"559" => q <= x"00";
            when x"55A" => q <= x"00";
            when x"55B" => q <= x"00";
            when x"55C" => q <= x"00";
            when x"55D" => q <= x"00";
            when x"55E" => q <= x"00";
            when x"55F" => q <= x"00";
            when x"560" => q <= x"00";
            when x"561" => q <= x"11";
            when x"562" => q <= x"11";
            when x"563" => q <= x"11";
            when x"564" => q <= x"0A";
            when x"565" => q <= x"0A";
            when x"566" => q <= x"04";
            when x"567" => q <= x"04";
            when x"568" => q <= x"00";
            when x"569" => q <= x"00";
            when x"56A" => q <= x"00";
            when x"56B" => q <= x"00";
            when x"56C" => q <= x"00";
            when x"56D" => q <= x"00";
            when x"56E" => q <= x"00";
            when x"56F" => q <= x"00";
            when x"570" => q <= x"00";
            when x"571" => q <= x"11";
            when x"572" => q <= x"11";
            when x"573" => q <= x"11";
            when x"574" => q <= x"15";
            when x"575" => q <= x"15";
            when x"576" => q <= x"15";
            when x"577" => q <= x"0A";
            when x"578" => q <= x"00";
            when x"579" => q <= x"00";
            when x"57A" => q <= x"00";
            when x"57B" => q <= x"00";
            when x"57C" => q <= x"00";
            when x"57D" => q <= x"00";
            when x"57E" => q <= x"00";
            when x"57F" => q <= x"00";
            when x"580" => q <= x"00";
            when x"581" => q <= x"11";
            when x"582" => q <= x"11";
            when x"583" => q <= x"0A";
            when x"584" => q <= x"04";
            when x"585" => q <= x"0A";
            when x"586" => q <= x"11";
            when x"587" => q <= x"11";
            when x"588" => q <= x"00";
            when x"589" => q <= x"00";
            when x"58A" => q <= x"00";
            when x"58B" => q <= x"00";
            when x"58C" => q <= x"00";
            when x"58D" => q <= x"00";
            when x"58E" => q <= x"00";
            when x"58F" => q <= x"00";
            when x"590" => q <= x"00";
            when x"591" => q <= x"11";
            when x"592" => q <= x"11";
            when x"593" => q <= x"0A";
            when x"594" => q <= x"04";
            when x"595" => q <= x"04";
            when x"596" => q <= x"04";
            when x"597" => q <= x"04";
            when x"598" => q <= x"00";
            when x"599" => q <= x"00";
            when x"59A" => q <= x"00";
            when x"59B" => q <= x"00";
            when x"59C" => q <= x"00";
            when x"59D" => q <= x"00";
            when x"59E" => q <= x"00";
            when x"59F" => q <= x"00";
            when x"5A0" => q <= x"00";
            when x"5A1" => q <= x"1F";
            when x"5A2" => q <= x"01";
            when x"5A3" => q <= x"02";
            when x"5A4" => q <= x"04";
            when x"5A5" => q <= x"08";
            when x"5A6" => q <= x"10";
            when x"5A7" => q <= x"1F";
            when x"5A8" => q <= x"00";
            when x"5A9" => q <= x"00";
            when x"5AA" => q <= x"00";
            when x"5AB" => q <= x"00";
            when x"5AC" => q <= x"00";
            when x"5AD" => q <= x"00";
            when x"5AE" => q <= x"00";
            when x"5AF" => q <= x"00";
            when x"5B0" => q <= x"00";
            when x"5B1" => q <= x"00";
            when x"5B2" => q <= x"04";
            when x"5B3" => q <= x"08";
            when x"5B4" => q <= x"1F";
            when x"5B5" => q <= x"08";
            when x"5B6" => q <= x"04";
            when x"5B7" => q <= x"00";
            when x"5B8" => q <= x"00";
            when x"5B9" => q <= x"00";
            when x"5BA" => q <= x"00";
            when x"5BB" => q <= x"00";
            when x"5BC" => q <= x"00";
            when x"5BD" => q <= x"00";
            when x"5BE" => q <= x"00";
            when x"5BF" => q <= x"00";
            when x"5C0" => q <= x"00";
            when x"5C1" => q <= x"10";
            when x"5C2" => q <= x"10";
            when x"5C3" => q <= x"10";
            when x"5C4" => q <= x"10";
            when x"5C5" => q <= x"16";
            when x"5C6" => q <= x"01";
            when x"5C7" => q <= x"02";
            when x"5C8" => q <= x"04";
            when x"5C9" => q <= x"07";
            when x"5CA" => q <= x"00";
            when x"5CB" => q <= x"00";
            when x"5CC" => q <= x"00";
            when x"5CD" => q <= x"00";
            when x"5CE" => q <= x"00";
            when x"5CF" => q <= x"00";
            when x"5D0" => q <= x"00";
            when x"5D1" => q <= x"00";
            when x"5D2" => q <= x"04";
            when x"5D3" => q <= x"02";
            when x"5D4" => q <= x"1F";
            when x"5D5" => q <= x"02";
            when x"5D6" => q <= x"04";
            when x"5D7" => q <= x"00";
            when x"5D8" => q <= x"00";
            when x"5D9" => q <= x"00";
            when x"5DA" => q <= x"00";
            when x"5DB" => q <= x"00";
            when x"5DC" => q <= x"00";
            when x"5DD" => q <= x"00";
            when x"5DE" => q <= x"00";
            when x"5DF" => q <= x"00";
            when x"5E0" => q <= x"00";
            when x"5E1" => q <= x"00";
            when x"5E2" => q <= x"04";
            when x"5E3" => q <= x"0E";
            when x"5E4" => q <= x"15";
            when x"5E5" => q <= x"04";
            when x"5E6" => q <= x"04";
            when x"5E7" => q <= x"00";
            when x"5E8" => q <= x"00";
            when x"5E9" => q <= x"00";
            when x"5EA" => q <= x"00";
            when x"5EB" => q <= x"00";
            when x"5EC" => q <= x"00";
            when x"5ED" => q <= x"00";
            when x"5EE" => q <= x"00";
            when x"5EF" => q <= x"00";
            when x"5F0" => q <= x"00";
            when x"5F1" => q <= x"0A";
            when x"5F2" => q <= x"0A";
            when x"5F3" => q <= x"1F";
            when x"5F4" => q <= x"0A";
            when x"5F5" => q <= x"1F";
            when x"5F6" => q <= x"0A";
            when x"5F7" => q <= x"0A";
            when x"5F8" => q <= x"00";
            when x"5F9" => q <= x"00";
            when x"5FA" => q <= x"00";
            when x"5FB" => q <= x"00";
            when x"5FC" => q <= x"00";
            when x"5FD" => q <= x"00";
            when x"5FE" => q <= x"00";
            when x"5FF" => q <= x"00";
            when x"600" => q <= x"00";
            when x"601" => q <= x"00";
            when x"602" => q <= x"00";
            when x"603" => q <= x"00";
            when x"604" => q <= x"1F";
            when x"605" => q <= x"00";
            when x"606" => q <= x"00";
            when x"607" => q <= x"00";
            when x"608" => q <= x"00";
            when x"609" => q <= x"00";
            when x"60A" => q <= x"00";
            when x"60B" => q <= x"00";
            when x"60C" => q <= x"00";
            when x"60D" => q <= x"00";
            when x"60E" => q <= x"00";
            when x"60F" => q <= x"00";
            when x"610" => q <= x"00";
            when x"611" => q <= x"00";
            when x"612" => q <= x"00";
            when x"613" => q <= x"0E";
            when x"614" => q <= x"01";
            when x"615" => q <= x"0F";
            when x"616" => q <= x"11";
            when x"617" => q <= x"0F";
            when x"618" => q <= x"00";
            when x"619" => q <= x"00";
            when x"61A" => q <= x"00";
            when x"61B" => q <= x"00";
            when x"61C" => q <= x"00";
            when x"61D" => q <= x"00";
            when x"61E" => q <= x"00";
            when x"61F" => q <= x"00";
            when x"620" => q <= x"00";
            when x"621" => q <= x"10";
            when x"622" => q <= x"10";
            when x"623" => q <= x"1E";
            when x"624" => q <= x"11";
            when x"625" => q <= x"11";
            when x"626" => q <= x"11";
            when x"627" => q <= x"1E";
            when x"628" => q <= x"00";
            when x"629" => q <= x"00";
            when x"62A" => q <= x"00";
            when x"62B" => q <= x"00";
            when x"62C" => q <= x"00";
            when x"62D" => q <= x"00";
            when x"62E" => q <= x"00";
            when x"62F" => q <= x"00";
            when x"630" => q <= x"00";
            when x"631" => q <= x"00";
            when x"632" => q <= x"00";
            when x"633" => q <= x"0F";
            when x"634" => q <= x"10";
            when x"635" => q <= x"10";
            when x"636" => q <= x"10";
            when x"637" => q <= x"0F";
            when x"638" => q <= x"00";
            when x"639" => q <= x"00";
            when x"63A" => q <= x"00";
            when x"63B" => q <= x"00";
            when x"63C" => q <= x"00";
            when x"63D" => q <= x"00";
            when x"63E" => q <= x"00";
            when x"63F" => q <= x"00";
            when x"640" => q <= x"00";
            when x"641" => q <= x"01";
            when x"642" => q <= x"01";
            when x"643" => q <= x"0F";
            when x"644" => q <= x"11";
            when x"645" => q <= x"11";
            when x"646" => q <= x"11";
            when x"647" => q <= x"0F";
            when x"648" => q <= x"00";
            when x"649" => q <= x"00";
            when x"64A" => q <= x"00";
            when x"64B" => q <= x"00";
            when x"64C" => q <= x"00";
            when x"64D" => q <= x"00";
            when x"64E" => q <= x"00";
            when x"64F" => q <= x"00";
            when x"650" => q <= x"00";
            when x"651" => q <= x"00";
            when x"652" => q <= x"00";
            when x"653" => q <= x"0E";
            when x"654" => q <= x"11";
            when x"655" => q <= x"1F";
            when x"656" => q <= x"10";
            when x"657" => q <= x"0E";
            when x"658" => q <= x"00";
            when x"659" => q <= x"00";
            when x"65A" => q <= x"00";
            when x"65B" => q <= x"00";
            when x"65C" => q <= x"00";
            when x"65D" => q <= x"00";
            when x"65E" => q <= x"00";
            when x"65F" => q <= x"00";
            when x"660" => q <= x"00";
            when x"661" => q <= x"02";
            when x"662" => q <= x"04";
            when x"663" => q <= x"04";
            when x"664" => q <= x"0E";
            when x"665" => q <= x"04";
            when x"666" => q <= x"04";
            when x"667" => q <= x"04";
            when x"668" => q <= x"00";
            when x"669" => q <= x"00";
            when x"66A" => q <= x"00";
            when x"66B" => q <= x"00";
            when x"66C" => q <= x"00";
            when x"66D" => q <= x"00";
            when x"66E" => q <= x"00";
            when x"66F" => q <= x"00";
            when x"670" => q <= x"00";
            when x"671" => q <= x"00";
            when x"672" => q <= x"00";
            when x"673" => q <= x"0F";
            when x"674" => q <= x"11";
            when x"675" => q <= x"11";
            when x"676" => q <= x"11";
            when x"677" => q <= x"0F";
            when x"678" => q <= x"01";
            when x"679" => q <= x"0E";
            when x"67A" => q <= x"00";
            when x"67B" => q <= x"00";
            when x"67C" => q <= x"00";
            when x"67D" => q <= x"00";
            when x"67E" => q <= x"00";
            when x"67F" => q <= x"00";
            when x"680" => q <= x"00";
            when x"681" => q <= x"10";
            when x"682" => q <= x"10";
            when x"683" => q <= x"1E";
            when x"684" => q <= x"11";
            when x"685" => q <= x"11";
            when x"686" => q <= x"11";
            when x"687" => q <= x"11";
            when x"688" => q <= x"00";
            when x"689" => q <= x"00";
            when x"68A" => q <= x"00";
            when x"68B" => q <= x"00";
            when x"68C" => q <= x"00";
            when x"68D" => q <= x"00";
            when x"68E" => q <= x"00";
            when x"68F" => q <= x"00";
            when x"690" => q <= x"00";
            when x"691" => q <= x"04";
            when x"692" => q <= x"00";
            when x"693" => q <= x"0C";
            when x"694" => q <= x"04";
            when x"695" => q <= x"04";
            when x"696" => q <= x"04";
            when x"697" => q <= x"0E";
            when x"698" => q <= x"00";
            when x"699" => q <= x"00";
            when x"69A" => q <= x"00";
            when x"69B" => q <= x"00";
            when x"69C" => q <= x"00";
            when x"69D" => q <= x"00";
            when x"69E" => q <= x"00";
            when x"69F" => q <= x"00";
            when x"6A0" => q <= x"00";
            when x"6A1" => q <= x"04";
            when x"6A2" => q <= x"00";
            when x"6A3" => q <= x"04";
            when x"6A4" => q <= x"04";
            when x"6A5" => q <= x"04";
            when x"6A6" => q <= x"04";
            when x"6A7" => q <= x"04";
            when x"6A8" => q <= x"04";
            when x"6A9" => q <= x"08";
            when x"6AA" => q <= x"00";
            when x"6AB" => q <= x"00";
            when x"6AC" => q <= x"00";
            when x"6AD" => q <= x"00";
            when x"6AE" => q <= x"00";
            when x"6AF" => q <= x"00";
            when x"6B0" => q <= x"00";
            when x"6B1" => q <= x"08";
            when x"6B2" => q <= x"08";
            when x"6B3" => q <= x"09";
            when x"6B4" => q <= x"0A";
            when x"6B5" => q <= x"0C";
            when x"6B6" => q <= x"0A";
            when x"6B7" => q <= x"09";
            when x"6B8" => q <= x"00";
            when x"6B9" => q <= x"00";
            when x"6BA" => q <= x"00";
            when x"6BB" => q <= x"00";
            when x"6BC" => q <= x"00";
            when x"6BD" => q <= x"00";
            when x"6BE" => q <= x"00";
            when x"6BF" => q <= x"00";
            when x"6C0" => q <= x"00";
            when x"6C1" => q <= x"0C";
            when x"6C2" => q <= x"04";
            when x"6C3" => q <= x"04";
            when x"6C4" => q <= x"04";
            when x"6C5" => q <= x"04";
            when x"6C6" => q <= x"04";
            when x"6C7" => q <= x"0E";
            when x"6C8" => q <= x"00";
            when x"6C9" => q <= x"00";
            when x"6CA" => q <= x"00";
            when x"6CB" => q <= x"00";
            when x"6CC" => q <= x"00";
            when x"6CD" => q <= x"00";
            when x"6CE" => q <= x"00";
            when x"6CF" => q <= x"00";
            when x"6D0" => q <= x"00";
            when x"6D1" => q <= x"00";
            when x"6D2" => q <= x"00";
            when x"6D3" => q <= x"1A";
            when x"6D4" => q <= x"15";
            when x"6D5" => q <= x"15";
            when x"6D6" => q <= x"15";
            when x"6D7" => q <= x"15";
            when x"6D8" => q <= x"00";
            when x"6D9" => q <= x"00";
            when x"6DA" => q <= x"00";
            when x"6DB" => q <= x"00";
            when x"6DC" => q <= x"00";
            when x"6DD" => q <= x"00";
            when x"6DE" => q <= x"00";
            when x"6DF" => q <= x"00";
            when x"6E0" => q <= x"00";
            when x"6E1" => q <= x"00";
            when x"6E2" => q <= x"00";
            when x"6E3" => q <= x"1E";
            when x"6E4" => q <= x"11";
            when x"6E5" => q <= x"11";
            when x"6E6" => q <= x"11";
            when x"6E7" => q <= x"11";
            when x"6E8" => q <= x"00";
            when x"6E9" => q <= x"00";
            when x"6EA" => q <= x"00";
            when x"6EB" => q <= x"00";
            when x"6EC" => q <= x"00";
            when x"6ED" => q <= x"00";
            when x"6EE" => q <= x"00";
            when x"6EF" => q <= x"00";
            when x"6F0" => q <= x"00";
            when x"6F1" => q <= x"00";
            when x"6F2" => q <= x"00";
            when x"6F3" => q <= x"0E";
            when x"6F4" => q <= x"11";
            when x"6F5" => q <= x"11";
            when x"6F6" => q <= x"11";
            when x"6F7" => q <= x"0E";
            when x"6F8" => q <= x"00";
            when x"6F9" => q <= x"00";
            when x"6FA" => q <= x"00";
            when x"6FB" => q <= x"00";
            when x"6FC" => q <= x"00";
            when x"6FD" => q <= x"00";
            when x"6FE" => q <= x"00";
            when x"6FF" => q <= x"00";
            when x"700" => q <= x"00";
            when x"701" => q <= x"00";
            when x"702" => q <= x"00";
            when x"703" => q <= x"1E";
            when x"704" => q <= x"11";
            when x"705" => q <= x"11";
            when x"706" => q <= x"11";
            when x"707" => q <= x"1E";
            when x"708" => q <= x"10";
            when x"709" => q <= x"10";
            when x"70A" => q <= x"00";
            when x"70B" => q <= x"00";
            when x"70C" => q <= x"00";
            when x"70D" => q <= x"00";
            when x"70E" => q <= x"00";
            when x"70F" => q <= x"00";
            when x"710" => q <= x"00";
            when x"711" => q <= x"00";
            when x"712" => q <= x"00";
            when x"713" => q <= x"0F";
            when x"714" => q <= x"11";
            when x"715" => q <= x"11";
            when x"716" => q <= x"11";
            when x"717" => q <= x"0F";
            when x"718" => q <= x"01";
            when x"719" => q <= x"01";
            when x"71A" => q <= x"00";
            when x"71B" => q <= x"00";
            when x"71C" => q <= x"00";
            when x"71D" => q <= x"00";
            when x"71E" => q <= x"00";
            when x"71F" => q <= x"00";
            when x"720" => q <= x"00";
            when x"721" => q <= x"00";
            when x"722" => q <= x"00";
            when x"723" => q <= x"0B";
            when x"724" => q <= x"0C";
            when x"725" => q <= x"08";
            when x"726" => q <= x"08";
            when x"727" => q <= x"08";
            when x"728" => q <= x"00";
            when x"729" => q <= x"00";
            when x"72A" => q <= x"00";
            when x"72B" => q <= x"00";
            when x"72C" => q <= x"00";
            when x"72D" => q <= x"00";
            when x"72E" => q <= x"00";
            when x"72F" => q <= x"00";
            when x"730" => q <= x"00";
            when x"731" => q <= x"00";
            when x"732" => q <= x"00";
            when x"733" => q <= x"0F";
            when x"734" => q <= x"10";
            when x"735" => q <= x"0E";
            when x"736" => q <= x"01";
            when x"737" => q <= x"1E";
            when x"738" => q <= x"00";
            when x"739" => q <= x"00";
            when x"73A" => q <= x"00";
            when x"73B" => q <= x"00";
            when x"73C" => q <= x"00";
            when x"73D" => q <= x"00";
            when x"73E" => q <= x"00";
            when x"73F" => q <= x"00";
            when x"740" => q <= x"00";
            when x"741" => q <= x"04";
            when x"742" => q <= x"04";
            when x"743" => q <= x"0E";
            when x"744" => q <= x"04";
            when x"745" => q <= x"04";
            when x"746" => q <= x"04";
            when x"747" => q <= x"02";
            when x"748" => q <= x"00";
            when x"749" => q <= x"00";
            when x"74A" => q <= x"00";
            when x"74B" => q <= x"00";
            when x"74C" => q <= x"00";
            when x"74D" => q <= x"00";
            when x"74E" => q <= x"00";
            when x"74F" => q <= x"00";
            when x"750" => q <= x"00";
            when x"751" => q <= x"00";
            when x"752" => q <= x"00";
            when x"753" => q <= x"11";
            when x"754" => q <= x"11";
            when x"755" => q <= x"11";
            when x"756" => q <= x"11";
            when x"757" => q <= x"0F";
            when x"758" => q <= x"00";
            when x"759" => q <= x"00";
            when x"75A" => q <= x"00";
            when x"75B" => q <= x"00";
            when x"75C" => q <= x"00";
            when x"75D" => q <= x"00";
            when x"75E" => q <= x"00";
            when x"75F" => q <= x"00";
            when x"760" => q <= x"00";
            when x"761" => q <= x"00";
            when x"762" => q <= x"00";
            when x"763" => q <= x"11";
            when x"764" => q <= x"11";
            when x"765" => q <= x"0A";
            when x"766" => q <= x"0A";
            when x"767" => q <= x"04";
            when x"768" => q <= x"00";
            when x"769" => q <= x"00";
            when x"76A" => q <= x"00";
            when x"76B" => q <= x"00";
            when x"76C" => q <= x"00";
            when x"76D" => q <= x"00";
            when x"76E" => q <= x"00";
            when x"76F" => q <= x"00";
            when x"770" => q <= x"00";
            when x"771" => q <= x"00";
            when x"772" => q <= x"00";
            when x"773" => q <= x"11";
            when x"774" => q <= x"11";
            when x"775" => q <= x"15";
            when x"776" => q <= x"15";
            when x"777" => q <= x"0A";
            when x"778" => q <= x"00";
            when x"779" => q <= x"00";
            when x"77A" => q <= x"00";
            when x"77B" => q <= x"00";
            when x"77C" => q <= x"00";
            when x"77D" => q <= x"00";
            when x"77E" => q <= x"00";
            when x"77F" => q <= x"00";
            when x"780" => q <= x"00";
            when x"781" => q <= x"00";
            when x"782" => q <= x"00";
            when x"783" => q <= x"11";
            when x"784" => q <= x"0A";
            when x"785" => q <= x"04";
            when x"786" => q <= x"0A";
            when x"787" => q <= x"11";
            when x"788" => q <= x"00";
            when x"789" => q <= x"00";
            when x"78A" => q <= x"00";
            when x"78B" => q <= x"00";
            when x"78C" => q <= x"00";
            when x"78D" => q <= x"00";
            when x"78E" => q <= x"00";
            when x"78F" => q <= x"00";
            when x"790" => q <= x"00";
            when x"791" => q <= x"00";
            when x"792" => q <= x"00";
            when x"793" => q <= x"11";
            when x"794" => q <= x"11";
            when x"795" => q <= x"11";
            when x"796" => q <= x"11";
            when x"797" => q <= x"0F";
            when x"798" => q <= x"01";
            when x"799" => q <= x"0E";
            when x"79A" => q <= x"00";
            when x"79B" => q <= x"00";
            when x"79C" => q <= x"00";
            when x"79D" => q <= x"00";
            when x"79E" => q <= x"00";
            when x"79F" => q <= x"00";
            when x"7A0" => q <= x"00";
            when x"7A1" => q <= x"00";
            when x"7A2" => q <= x"00";
            when x"7A3" => q <= x"1F";
            when x"7A4" => q <= x"02";
            when x"7A5" => q <= x"04";
            when x"7A6" => q <= x"08";
            when x"7A7" => q <= x"1F";
            when x"7A8" => q <= x"00";
            when x"7A9" => q <= x"00";
            when x"7AA" => q <= x"00";
            when x"7AB" => q <= x"00";
            when x"7AC" => q <= x"00";
            when x"7AD" => q <= x"00";
            when x"7AE" => q <= x"00";
            when x"7AF" => q <= x"00";
            when x"7B0" => q <= x"00";
            when x"7B1" => q <= x"08";
            when x"7B2" => q <= x"08";
            when x"7B3" => q <= x"08";
            when x"7B4" => q <= x"08";
            when x"7B5" => q <= x"09";
            when x"7B6" => q <= x"03";
            when x"7B7" => q <= x"05";
            when x"7B8" => q <= x"07";
            when x"7B9" => q <= x"01";
            when x"7BA" => q <= x"00";
            when x"7BB" => q <= x"00";
            when x"7BC" => q <= x"00";
            when x"7BD" => q <= x"00";
            when x"7BE" => q <= x"00";
            when x"7BF" => q <= x"00";
            when x"7C0" => q <= x"00";
            when x"7C1" => q <= x"0A";
            when x"7C2" => q <= x"0A";
            when x"7C3" => q <= x"0A";
            when x"7C4" => q <= x"0A";
            when x"7C5" => q <= x"0A";
            when x"7C6" => q <= x"0A";
            when x"7C7" => q <= x"0A";
            when x"7C8" => q <= x"00";
            when x"7C9" => q <= x"00";
            when x"7CA" => q <= x"00";
            when x"7CB" => q <= x"00";
            when x"7CC" => q <= x"00";
            when x"7CD" => q <= x"00";
            when x"7CE" => q <= x"00";
            when x"7CF" => q <= x"00";
            when x"7D0" => q <= x"00";
            when x"7D1" => q <= x"18";
            when x"7D2" => q <= x"04";
            when x"7D3" => q <= x"18";
            when x"7D4" => q <= x"04";
            when x"7D5" => q <= x"19";
            when x"7D6" => q <= x"03";
            when x"7D7" => q <= x"05";
            when x"7D8" => q <= x"07";
            when x"7D9" => q <= x"01";
            when x"7DA" => q <= x"00";
            when x"7DB" => q <= x"00";
            when x"7DC" => q <= x"00";
            when x"7DD" => q <= x"00";
            when x"7DE" => q <= x"00";
            when x"7DF" => q <= x"00";
            when x"7E0" => q <= x"00";
            when x"7E1" => q <= x"00";
            when x"7E2" => q <= x"04";
            when x"7E3" => q <= x"00";
            when x"7E4" => q <= x"1F";
            when x"7E5" => q <= x"00";
            when x"7E6" => q <= x"04";
            when x"7E7" => q <= x"00";
            when x"7E8" => q <= x"00";
            when x"7E9" => q <= x"00";
            when x"7EA" => q <= x"00";
            when x"7EB" => q <= x"00";
            when x"7EC" => q <= x"00";
            when x"7ED" => q <= x"00";
            when x"7EE" => q <= x"00";
            when x"7EF" => q <= x"00";
            when x"7F0" => q <= x"00";
            when x"7F1" => q <= x"1F";
            when x"7F2" => q <= x"1F";
            when x"7F3" => q <= x"1F";
            when x"7F4" => q <= x"1F";
            when x"7F5" => q <= x"1F";
            when x"7F6" => q <= x"1F";
            when x"7F7" => q <= x"1F";
            when x"7F8" => q <= x"00";
            when x"7F9" => q <= x"00";
            when x"7FA" => q <= x"00";
            when x"7FB" => q <= x"00";
            when x"7FC" => q <= x"00";
            when x"7FD" => q <= x"00";
            when x"7FE" => q <= x"00";
            when x"7FF" => q <= x"00";
            when x"800" => q <= x"00";
            when x"801" => q <= x"00";
            when x"802" => q <= x"00";
            when x"803" => q <= x"00";
            when x"804" => q <= x"00";
            when x"805" => q <= x"00";
            when x"806" => q <= x"00";
            when x"807" => q <= x"00";
            when x"808" => q <= x"00";
            when x"809" => q <= x"00";
            when x"80A" => q <= x"00";
            when x"80B" => q <= x"00";
            when x"80C" => q <= x"00";
            when x"80D" => q <= x"00";
            when x"80E" => q <= x"00";
            when x"80F" => q <= x"00";
            when x"810" => q <= x"00";
            when x"811" => q <= x"00";
            when x"812" => q <= x"00";
            when x"813" => q <= x"00";
            when x"814" => q <= x"00";
            when x"815" => q <= x"00";
            when x"816" => q <= x"00";
            when x"817" => q <= x"00";
            when x"818" => q <= x"00";
            when x"819" => q <= x"00";
            when x"81A" => q <= x"00";
            when x"81B" => q <= x"00";
            when x"81C" => q <= x"00";
            when x"81D" => q <= x"00";
            when x"81E" => q <= x"00";
            when x"81F" => q <= x"00";
            when x"820" => q <= x"00";
            when x"821" => q <= x"00";
            when x"822" => q <= x"00";
            when x"823" => q <= x"00";
            when x"824" => q <= x"00";
            when x"825" => q <= x"00";
            when x"826" => q <= x"00";
            when x"827" => q <= x"00";
            when x"828" => q <= x"00";
            when x"829" => q <= x"00";
            when x"82A" => q <= x"00";
            when x"82B" => q <= x"00";
            when x"82C" => q <= x"00";
            when x"82D" => q <= x"00";
            when x"82E" => q <= x"00";
            when x"82F" => q <= x"00";
            when x"830" => q <= x"00";
            when x"831" => q <= x"00";
            when x"832" => q <= x"00";
            when x"833" => q <= x"00";
            when x"834" => q <= x"00";
            when x"835" => q <= x"00";
            when x"836" => q <= x"00";
            when x"837" => q <= x"00";
            when x"838" => q <= x"00";
            when x"839" => q <= x"00";
            when x"83A" => q <= x"00";
            when x"83B" => q <= x"00";
            when x"83C" => q <= x"00";
            when x"83D" => q <= x"00";
            when x"83E" => q <= x"00";
            when x"83F" => q <= x"00";
            when x"840" => q <= x"00";
            when x"841" => q <= x"00";
            when x"842" => q <= x"00";
            when x"843" => q <= x"00";
            when x"844" => q <= x"00";
            when x"845" => q <= x"00";
            when x"846" => q <= x"00";
            when x"847" => q <= x"00";
            when x"848" => q <= x"00";
            when x"849" => q <= x"00";
            when x"84A" => q <= x"00";
            when x"84B" => q <= x"00";
            when x"84C" => q <= x"00";
            when x"84D" => q <= x"00";
            when x"84E" => q <= x"00";
            when x"84F" => q <= x"00";
            when x"850" => q <= x"00";
            when x"851" => q <= x"00";
            when x"852" => q <= x"00";
            when x"853" => q <= x"00";
            when x"854" => q <= x"00";
            when x"855" => q <= x"00";
            when x"856" => q <= x"00";
            when x"857" => q <= x"00";
            when x"858" => q <= x"00";
            when x"859" => q <= x"00";
            when x"85A" => q <= x"00";
            when x"85B" => q <= x"00";
            when x"85C" => q <= x"00";
            when x"85D" => q <= x"00";
            when x"85E" => q <= x"00";
            when x"85F" => q <= x"00";
            when x"860" => q <= x"00";
            when x"861" => q <= x"00";
            when x"862" => q <= x"00";
            when x"863" => q <= x"00";
            when x"864" => q <= x"00";
            when x"865" => q <= x"00";
            when x"866" => q <= x"00";
            when x"867" => q <= x"00";
            when x"868" => q <= x"00";
            when x"869" => q <= x"00";
            when x"86A" => q <= x"00";
            when x"86B" => q <= x"00";
            when x"86C" => q <= x"00";
            when x"86D" => q <= x"00";
            when x"86E" => q <= x"00";
            when x"86F" => q <= x"00";
            when x"870" => q <= x"00";
            when x"871" => q <= x"00";
            when x"872" => q <= x"00";
            when x"873" => q <= x"00";
            when x"874" => q <= x"00";
            when x"875" => q <= x"00";
            when x"876" => q <= x"00";
            when x"877" => q <= x"00";
            when x"878" => q <= x"00";
            when x"879" => q <= x"00";
            when x"87A" => q <= x"00";
            when x"87B" => q <= x"00";
            when x"87C" => q <= x"00";
            when x"87D" => q <= x"00";
            when x"87E" => q <= x"00";
            when x"87F" => q <= x"00";
            when x"880" => q <= x"00";
            when x"881" => q <= x"00";
            when x"882" => q <= x"00";
            when x"883" => q <= x"00";
            when x"884" => q <= x"00";
            when x"885" => q <= x"00";
            when x"886" => q <= x"00";
            when x"887" => q <= x"00";
            when x"888" => q <= x"00";
            when x"889" => q <= x"00";
            when x"88A" => q <= x"00";
            when x"88B" => q <= x"00";
            when x"88C" => q <= x"00";
            when x"88D" => q <= x"00";
            when x"88E" => q <= x"00";
            when x"88F" => q <= x"00";
            when x"890" => q <= x"00";
            when x"891" => q <= x"00";
            when x"892" => q <= x"00";
            when x"893" => q <= x"00";
            when x"894" => q <= x"00";
            when x"895" => q <= x"00";
            when x"896" => q <= x"00";
            when x"897" => q <= x"00";
            when x"898" => q <= x"00";
            when x"899" => q <= x"00";
            when x"89A" => q <= x"00";
            when x"89B" => q <= x"00";
            when x"89C" => q <= x"00";
            when x"89D" => q <= x"00";
            when x"89E" => q <= x"00";
            when x"89F" => q <= x"00";
            when x"8A0" => q <= x"00";
            when x"8A1" => q <= x"00";
            when x"8A2" => q <= x"00";
            when x"8A3" => q <= x"00";
            when x"8A4" => q <= x"00";
            when x"8A5" => q <= x"00";
            when x"8A6" => q <= x"00";
            when x"8A7" => q <= x"00";
            when x"8A8" => q <= x"00";
            when x"8A9" => q <= x"00";
            when x"8AA" => q <= x"00";
            when x"8AB" => q <= x"00";
            when x"8AC" => q <= x"00";
            when x"8AD" => q <= x"00";
            when x"8AE" => q <= x"00";
            when x"8AF" => q <= x"00";
            when x"8B0" => q <= x"00";
            when x"8B1" => q <= x"00";
            when x"8B2" => q <= x"00";
            when x"8B3" => q <= x"00";
            when x"8B4" => q <= x"00";
            when x"8B5" => q <= x"00";
            when x"8B6" => q <= x"00";
            when x"8B7" => q <= x"00";
            when x"8B8" => q <= x"00";
            when x"8B9" => q <= x"00";
            when x"8BA" => q <= x"00";
            when x"8BB" => q <= x"00";
            when x"8BC" => q <= x"00";
            when x"8BD" => q <= x"00";
            when x"8BE" => q <= x"00";
            when x"8BF" => q <= x"00";
            when x"8C0" => q <= x"00";
            when x"8C1" => q <= x"00";
            when x"8C2" => q <= x"00";
            when x"8C3" => q <= x"00";
            when x"8C4" => q <= x"00";
            when x"8C5" => q <= x"00";
            when x"8C6" => q <= x"00";
            when x"8C7" => q <= x"00";
            when x"8C8" => q <= x"00";
            when x"8C9" => q <= x"00";
            when x"8CA" => q <= x"00";
            when x"8CB" => q <= x"00";
            when x"8CC" => q <= x"00";
            when x"8CD" => q <= x"00";
            when x"8CE" => q <= x"00";
            when x"8CF" => q <= x"00";
            when x"8D0" => q <= x"00";
            when x"8D1" => q <= x"00";
            when x"8D2" => q <= x"00";
            when x"8D3" => q <= x"00";
            when x"8D4" => q <= x"00";
            when x"8D5" => q <= x"00";
            when x"8D6" => q <= x"00";
            when x"8D7" => q <= x"00";
            when x"8D8" => q <= x"00";
            when x"8D9" => q <= x"00";
            when x"8DA" => q <= x"00";
            when x"8DB" => q <= x"00";
            when x"8DC" => q <= x"00";
            when x"8DD" => q <= x"00";
            when x"8DE" => q <= x"00";
            when x"8DF" => q <= x"00";
            when x"8E0" => q <= x"00";
            when x"8E1" => q <= x"00";
            when x"8E2" => q <= x"00";
            when x"8E3" => q <= x"00";
            when x"8E4" => q <= x"00";
            when x"8E5" => q <= x"00";
            when x"8E6" => q <= x"00";
            when x"8E7" => q <= x"00";
            when x"8E8" => q <= x"00";
            when x"8E9" => q <= x"00";
            when x"8EA" => q <= x"00";
            when x"8EB" => q <= x"00";
            when x"8EC" => q <= x"00";
            when x"8ED" => q <= x"00";
            when x"8EE" => q <= x"00";
            when x"8EF" => q <= x"00";
            when x"8F0" => q <= x"00";
            when x"8F1" => q <= x"00";
            when x"8F2" => q <= x"00";
            when x"8F3" => q <= x"00";
            when x"8F4" => q <= x"00";
            when x"8F5" => q <= x"00";
            when x"8F6" => q <= x"00";
            when x"8F7" => q <= x"00";
            when x"8F8" => q <= x"00";
            when x"8F9" => q <= x"00";
            when x"8FA" => q <= x"00";
            when x"8FB" => q <= x"00";
            when x"8FC" => q <= x"00";
            when x"8FD" => q <= x"00";
            when x"8FE" => q <= x"00";
            when x"8FF" => q <= x"00";
            when x"900" => q <= x"00";
            when x"901" => q <= x"00";
            when x"902" => q <= x"00";
            when x"903" => q <= x"00";
            when x"904" => q <= x"00";
            when x"905" => q <= x"00";
            when x"906" => q <= x"00";
            when x"907" => q <= x"00";
            when x"908" => q <= x"00";
            when x"909" => q <= x"00";
            when x"90A" => q <= x"00";
            when x"90B" => q <= x"00";
            when x"90C" => q <= x"00";
            when x"90D" => q <= x"00";
            when x"90E" => q <= x"00";
            when x"90F" => q <= x"00";
            when x"910" => q <= x"00";
            when x"911" => q <= x"00";
            when x"912" => q <= x"00";
            when x"913" => q <= x"00";
            when x"914" => q <= x"00";
            when x"915" => q <= x"00";
            when x"916" => q <= x"00";
            when x"917" => q <= x"00";
            when x"918" => q <= x"00";
            when x"919" => q <= x"00";
            when x"91A" => q <= x"00";
            when x"91B" => q <= x"00";
            when x"91C" => q <= x"00";
            when x"91D" => q <= x"00";
            when x"91E" => q <= x"00";
            when x"91F" => q <= x"00";
            when x"920" => q <= x"00";
            when x"921" => q <= x"00";
            when x"922" => q <= x"00";
            when x"923" => q <= x"00";
            when x"924" => q <= x"00";
            when x"925" => q <= x"00";
            when x"926" => q <= x"00";
            when x"927" => q <= x"00";
            when x"928" => q <= x"00";
            when x"929" => q <= x"00";
            when x"92A" => q <= x"00";
            when x"92B" => q <= x"00";
            when x"92C" => q <= x"00";
            when x"92D" => q <= x"00";
            when x"92E" => q <= x"00";
            when x"92F" => q <= x"00";
            when x"930" => q <= x"00";
            when x"931" => q <= x"00";
            when x"932" => q <= x"00";
            when x"933" => q <= x"00";
            when x"934" => q <= x"00";
            when x"935" => q <= x"00";
            when x"936" => q <= x"00";
            when x"937" => q <= x"00";
            when x"938" => q <= x"00";
            when x"939" => q <= x"00";
            when x"93A" => q <= x"00";
            when x"93B" => q <= x"00";
            when x"93C" => q <= x"00";
            when x"93D" => q <= x"00";
            when x"93E" => q <= x"00";
            when x"93F" => q <= x"00";
            when x"940" => q <= x"00";
            when x"941" => q <= x"00";
            when x"942" => q <= x"00";
            when x"943" => q <= x"00";
            when x"944" => q <= x"00";
            when x"945" => q <= x"00";
            when x"946" => q <= x"00";
            when x"947" => q <= x"00";
            when x"948" => q <= x"00";
            when x"949" => q <= x"00";
            when x"94A" => q <= x"00";
            when x"94B" => q <= x"00";
            when x"94C" => q <= x"00";
            when x"94D" => q <= x"00";
            when x"94E" => q <= x"00";
            when x"94F" => q <= x"00";
            when x"950" => q <= x"00";
            when x"951" => q <= x"00";
            when x"952" => q <= x"00";
            when x"953" => q <= x"00";
            when x"954" => q <= x"00";
            when x"955" => q <= x"00";
            when x"956" => q <= x"00";
            when x"957" => q <= x"00";
            when x"958" => q <= x"00";
            when x"959" => q <= x"00";
            when x"95A" => q <= x"00";
            when x"95B" => q <= x"00";
            when x"95C" => q <= x"00";
            when x"95D" => q <= x"00";
            when x"95E" => q <= x"00";
            when x"95F" => q <= x"00";
            when x"960" => q <= x"00";
            when x"961" => q <= x"00";
            when x"962" => q <= x"00";
            when x"963" => q <= x"00";
            when x"964" => q <= x"00";
            when x"965" => q <= x"00";
            when x"966" => q <= x"00";
            when x"967" => q <= x"00";
            when x"968" => q <= x"00";
            when x"969" => q <= x"00";
            when x"96A" => q <= x"00";
            when x"96B" => q <= x"00";
            when x"96C" => q <= x"00";
            when x"96D" => q <= x"00";
            when x"96E" => q <= x"00";
            when x"96F" => q <= x"00";
            when x"970" => q <= x"00";
            when x"971" => q <= x"00";
            when x"972" => q <= x"00";
            when x"973" => q <= x"00";
            when x"974" => q <= x"00";
            when x"975" => q <= x"00";
            when x"976" => q <= x"00";
            when x"977" => q <= x"00";
            when x"978" => q <= x"00";
            when x"979" => q <= x"00";
            when x"97A" => q <= x"00";
            when x"97B" => q <= x"00";
            when x"97C" => q <= x"00";
            when x"97D" => q <= x"00";
            when x"97E" => q <= x"00";
            when x"97F" => q <= x"00";
            when x"980" => q <= x"00";
            when x"981" => q <= x"00";
            when x"982" => q <= x"00";
            when x"983" => q <= x"00";
            when x"984" => q <= x"00";
            when x"985" => q <= x"00";
            when x"986" => q <= x"00";
            when x"987" => q <= x"00";
            when x"988" => q <= x"00";
            when x"989" => q <= x"00";
            when x"98A" => q <= x"00";
            when x"98B" => q <= x"00";
            when x"98C" => q <= x"00";
            when x"98D" => q <= x"00";
            when x"98E" => q <= x"00";
            when x"98F" => q <= x"00";
            when x"990" => q <= x"00";
            when x"991" => q <= x"00";
            when x"992" => q <= x"00";
            when x"993" => q <= x"00";
            when x"994" => q <= x"00";
            when x"995" => q <= x"00";
            when x"996" => q <= x"00";
            when x"997" => q <= x"00";
            when x"998" => q <= x"00";
            when x"999" => q <= x"00";
            when x"99A" => q <= x"00";
            when x"99B" => q <= x"00";
            when x"99C" => q <= x"00";
            when x"99D" => q <= x"00";
            when x"99E" => q <= x"00";
            when x"99F" => q <= x"00";
            when x"9A0" => q <= x"00";
            when x"9A1" => q <= x"00";
            when x"9A2" => q <= x"00";
            when x"9A3" => q <= x"00";
            when x"9A4" => q <= x"00";
            when x"9A5" => q <= x"00";
            when x"9A6" => q <= x"00";
            when x"9A7" => q <= x"00";
            when x"9A8" => q <= x"00";
            when x"9A9" => q <= x"00";
            when x"9AA" => q <= x"00";
            when x"9AB" => q <= x"00";
            when x"9AC" => q <= x"00";
            when x"9AD" => q <= x"00";
            when x"9AE" => q <= x"00";
            when x"9AF" => q <= x"00";
            when x"9B0" => q <= x"00";
            when x"9B1" => q <= x"00";
            when x"9B2" => q <= x"00";
            when x"9B3" => q <= x"00";
            when x"9B4" => q <= x"00";
            when x"9B5" => q <= x"00";
            when x"9B6" => q <= x"00";
            when x"9B7" => q <= x"00";
            when x"9B8" => q <= x"00";
            when x"9B9" => q <= x"00";
            when x"9BA" => q <= x"00";
            when x"9BB" => q <= x"00";
            when x"9BC" => q <= x"00";
            when x"9BD" => q <= x"00";
            when x"9BE" => q <= x"00";
            when x"9BF" => q <= x"00";
            when x"9C0" => q <= x"00";
            when x"9C1" => q <= x"00";
            when x"9C2" => q <= x"00";
            when x"9C3" => q <= x"00";
            when x"9C4" => q <= x"00";
            when x"9C5" => q <= x"00";
            when x"9C6" => q <= x"00";
            when x"9C7" => q <= x"00";
            when x"9C8" => q <= x"00";
            when x"9C9" => q <= x"00";
            when x"9CA" => q <= x"00";
            when x"9CB" => q <= x"00";
            when x"9CC" => q <= x"00";
            when x"9CD" => q <= x"00";
            when x"9CE" => q <= x"00";
            when x"9CF" => q <= x"00";
            when x"9D0" => q <= x"00";
            when x"9D1" => q <= x"00";
            when x"9D2" => q <= x"00";
            when x"9D3" => q <= x"00";
            when x"9D4" => q <= x"00";
            when x"9D5" => q <= x"00";
            when x"9D6" => q <= x"00";
            when x"9D7" => q <= x"00";
            when x"9D8" => q <= x"00";
            when x"9D9" => q <= x"00";
            when x"9DA" => q <= x"00";
            when x"9DB" => q <= x"00";
            when x"9DC" => q <= x"00";
            when x"9DD" => q <= x"00";
            when x"9DE" => q <= x"00";
            when x"9DF" => q <= x"00";
            when x"9E0" => q <= x"00";
            when x"9E1" => q <= x"00";
            when x"9E2" => q <= x"00";
            when x"9E3" => q <= x"00";
            when x"9E4" => q <= x"00";
            when x"9E5" => q <= x"00";
            when x"9E6" => q <= x"00";
            when x"9E7" => q <= x"00";
            when x"9E8" => q <= x"00";
            when x"9E9" => q <= x"00";
            when x"9EA" => q <= x"00";
            when x"9EB" => q <= x"00";
            when x"9EC" => q <= x"00";
            when x"9ED" => q <= x"00";
            when x"9EE" => q <= x"00";
            when x"9EF" => q <= x"00";
            when x"9F0" => q <= x"00";
            when x"9F1" => q <= x"00";
            when x"9F2" => q <= x"00";
            when x"9F3" => q <= x"00";
            when x"9F4" => q <= x"00";
            when x"9F5" => q <= x"00";
            when x"9F6" => q <= x"00";
            when x"9F7" => q <= x"00";
            when x"9F8" => q <= x"00";
            when x"9F9" => q <= x"00";
            when x"9FA" => q <= x"00";
            when x"9FB" => q <= x"00";
            when x"9FC" => q <= x"00";
            when x"9FD" => q <= x"00";
            when x"9FE" => q <= x"00";
            when x"9FF" => q <= x"00";
            when x"A00" => q <= x"80";
            when x"A01" => q <= x"80";
            when x"A02" => q <= x"80";
            when x"A03" => q <= x"80";
            when x"A04" => q <= x"80";
            when x"A05" => q <= x"80";
            when x"A06" => q <= x"80";
            when x"A07" => q <= x"80";
            when x"A08" => q <= x"80";
            when x"A09" => q <= x"80";
            when x"A0A" => q <= x"00";
            when x"A0B" => q <= x"00";
            when x"A0C" => q <= x"00";
            when x"A0D" => q <= x"00";
            when x"A0E" => q <= x"00";
            when x"A0F" => q <= x"00";
            when x"A10" => q <= x"B8";
            when x"A11" => q <= x"B8";
            when x"A12" => q <= x"B8";
            when x"A13" => q <= x"80";
            when x"A14" => q <= x"80";
            when x"A15" => q <= x"80";
            when x"A16" => q <= x"80";
            when x"A17" => q <= x"80";
            when x"A18" => q <= x"80";
            when x"A19" => q <= x"80";
            when x"A1A" => q <= x"00";
            when x"A1B" => q <= x"00";
            when x"A1C" => q <= x"00";
            when x"A1D" => q <= x"00";
            when x"A1E" => q <= x"00";
            when x"A1F" => q <= x"00";
            when x"A20" => q <= x"87";
            when x"A21" => q <= x"87";
            when x"A22" => q <= x"87";
            when x"A23" => q <= x"80";
            when x"A24" => q <= x"80";
            when x"A25" => q <= x"80";
            when x"A26" => q <= x"80";
            when x"A27" => q <= x"80";
            when x"A28" => q <= x"80";
            when x"A29" => q <= x"80";
            when x"A2A" => q <= x"00";
            when x"A2B" => q <= x"00";
            when x"A2C" => q <= x"00";
            when x"A2D" => q <= x"00";
            when x"A2E" => q <= x"00";
            when x"A2F" => q <= x"00";
            when x"A30" => q <= x"BF";
            when x"A31" => q <= x"BF";
            when x"A32" => q <= x"BF";
            when x"A33" => q <= x"80";
            when x"A34" => q <= x"80";
            when x"A35" => q <= x"80";
            when x"A36" => q <= x"80";
            when x"A37" => q <= x"80";
            when x"A38" => q <= x"80";
            when x"A39" => q <= x"80";
            when x"A3A" => q <= x"00";
            when x"A3B" => q <= x"00";
            when x"A3C" => q <= x"00";
            when x"A3D" => q <= x"00";
            when x"A3E" => q <= x"00";
            when x"A3F" => q <= x"00";
            when x"A40" => q <= x"80";
            when x"A41" => q <= x"80";
            when x"A42" => q <= x"80";
            when x"A43" => q <= x"B8";
            when x"A44" => q <= x"B8";
            when x"A45" => q <= x"B8";
            when x"A46" => q <= x"B8";
            when x"A47" => q <= x"80";
            when x"A48" => q <= x"80";
            when x"A49" => q <= x"80";
            when x"A4A" => q <= x"00";
            when x"A4B" => q <= x"00";
            when x"A4C" => q <= x"00";
            when x"A4D" => q <= x"00";
            when x"A4E" => q <= x"00";
            when x"A4F" => q <= x"00";
            when x"A50" => q <= x"B8";
            when x"A51" => q <= x"B8";
            when x"A52" => q <= x"B8";
            when x"A53" => q <= x"B8";
            when x"A54" => q <= x"B8";
            when x"A55" => q <= x"B8";
            when x"A56" => q <= x"B8";
            when x"A57" => q <= x"80";
            when x"A58" => q <= x"80";
            when x"A59" => q <= x"80";
            when x"A5A" => q <= x"00";
            when x"A5B" => q <= x"00";
            when x"A5C" => q <= x"00";
            when x"A5D" => q <= x"00";
            when x"A5E" => q <= x"00";
            when x"A5F" => q <= x"00";
            when x"A60" => q <= x"87";
            when x"A61" => q <= x"87";
            when x"A62" => q <= x"87";
            when x"A63" => q <= x"B8";
            when x"A64" => q <= x"B8";
            when x"A65" => q <= x"B8";
            when x"A66" => q <= x"B8";
            when x"A67" => q <= x"80";
            when x"A68" => q <= x"80";
            when x"A69" => q <= x"80";
            when x"A6A" => q <= x"00";
            when x"A6B" => q <= x"00";
            when x"A6C" => q <= x"00";
            when x"A6D" => q <= x"00";
            when x"A6E" => q <= x"00";
            when x"A6F" => q <= x"00";
            when x"A70" => q <= x"BF";
            when x"A71" => q <= x"BF";
            when x"A72" => q <= x"BF";
            when x"A73" => q <= x"B8";
            when x"A74" => q <= x"B8";
            when x"A75" => q <= x"B8";
            when x"A76" => q <= x"B8";
            when x"A77" => q <= x"80";
            when x"A78" => q <= x"80";
            when x"A79" => q <= x"80";
            when x"A7A" => q <= x"00";
            when x"A7B" => q <= x"00";
            when x"A7C" => q <= x"00";
            when x"A7D" => q <= x"00";
            when x"A7E" => q <= x"00";
            when x"A7F" => q <= x"00";
            when x"A80" => q <= x"80";
            when x"A81" => q <= x"80";
            when x"A82" => q <= x"80";
            when x"A83" => q <= x"87";
            when x"A84" => q <= x"87";
            when x"A85" => q <= x"87";
            when x"A86" => q <= x"87";
            when x"A87" => q <= x"80";
            when x"A88" => q <= x"80";
            when x"A89" => q <= x"80";
            when x"A8A" => q <= x"00";
            when x"A8B" => q <= x"00";
            when x"A8C" => q <= x"00";
            when x"A8D" => q <= x"00";
            when x"A8E" => q <= x"00";
            when x"A8F" => q <= x"00";
            when x"A90" => q <= x"B8";
            when x"A91" => q <= x"B8";
            when x"A92" => q <= x"B8";
            when x"A93" => q <= x"87";
            when x"A94" => q <= x"87";
            when x"A95" => q <= x"87";
            when x"A96" => q <= x"87";
            when x"A97" => q <= x"80";
            when x"A98" => q <= x"80";
            when x"A99" => q <= x"80";
            when x"A9A" => q <= x"00";
            when x"A9B" => q <= x"00";
            when x"A9C" => q <= x"00";
            when x"A9D" => q <= x"00";
            when x"A9E" => q <= x"00";
            when x"A9F" => q <= x"00";
            when x"AA0" => q <= x"87";
            when x"AA1" => q <= x"87";
            when x"AA2" => q <= x"87";
            when x"AA3" => q <= x"87";
            when x"AA4" => q <= x"87";
            when x"AA5" => q <= x"87";
            when x"AA6" => q <= x"87";
            when x"AA7" => q <= x"80";
            when x"AA8" => q <= x"80";
            when x"AA9" => q <= x"80";
            when x"AAA" => q <= x"00";
            when x"AAB" => q <= x"00";
            when x"AAC" => q <= x"00";
            when x"AAD" => q <= x"00";
            when x"AAE" => q <= x"00";
            when x"AAF" => q <= x"00";
            when x"AB0" => q <= x"BF";
            when x"AB1" => q <= x"BF";
            when x"AB2" => q <= x"BF";
            when x"AB3" => q <= x"87";
            when x"AB4" => q <= x"87";
            when x"AB5" => q <= x"87";
            when x"AB6" => q <= x"87";
            when x"AB7" => q <= x"80";
            when x"AB8" => q <= x"80";
            when x"AB9" => q <= x"80";
            when x"ABA" => q <= x"00";
            when x"ABB" => q <= x"00";
            when x"ABC" => q <= x"00";
            when x"ABD" => q <= x"00";
            when x"ABE" => q <= x"00";
            when x"ABF" => q <= x"00";
            when x"AC0" => q <= x"80";
            when x"AC1" => q <= x"80";
            when x"AC2" => q <= x"80";
            when x"AC3" => q <= x"BF";
            when x"AC4" => q <= x"BF";
            when x"AC5" => q <= x"BF";
            when x"AC6" => q <= x"BF";
            when x"AC7" => q <= x"80";
            when x"AC8" => q <= x"80";
            when x"AC9" => q <= x"80";
            when x"ACA" => q <= x"00";
            when x"ACB" => q <= x"00";
            when x"ACC" => q <= x"00";
            when x"ACD" => q <= x"00";
            when x"ACE" => q <= x"00";
            when x"ACF" => q <= x"00";
            when x"AD0" => q <= x"B8";
            when x"AD1" => q <= x"B8";
            when x"AD2" => q <= x"B8";
            when x"AD3" => q <= x"BF";
            when x"AD4" => q <= x"BF";
            when x"AD5" => q <= x"BF";
            when x"AD6" => q <= x"BF";
            when x"AD7" => q <= x"80";
            when x"AD8" => q <= x"80";
            when x"AD9" => q <= x"80";
            when x"ADA" => q <= x"00";
            when x"ADB" => q <= x"00";
            when x"ADC" => q <= x"00";
            when x"ADD" => q <= x"00";
            when x"ADE" => q <= x"00";
            when x"ADF" => q <= x"00";
            when x"AE0" => q <= x"87";
            when x"AE1" => q <= x"87";
            when x"AE2" => q <= x"87";
            when x"AE3" => q <= x"BF";
            when x"AE4" => q <= x"BF";
            when x"AE5" => q <= x"BF";
            when x"AE6" => q <= x"BF";
            when x"AE7" => q <= x"80";
            when x"AE8" => q <= x"80";
            when x"AE9" => q <= x"80";
            when x"AEA" => q <= x"00";
            when x"AEB" => q <= x"00";
            when x"AEC" => q <= x"00";
            when x"AED" => q <= x"00";
            when x"AEE" => q <= x"00";
            when x"AEF" => q <= x"00";
            when x"AF0" => q <= x"BF";
            when x"AF1" => q <= x"BF";
            when x"AF2" => q <= x"BF";
            when x"AF3" => q <= x"BF";
            when x"AF4" => q <= x"BF";
            when x"AF5" => q <= x"BF";
            when x"AF6" => q <= x"BF";
            when x"AF7" => q <= x"80";
            when x"AF8" => q <= x"80";
            when x"AF9" => q <= x"80";
            when x"AFA" => q <= x"00";
            when x"AFB" => q <= x"00";
            when x"AFC" => q <= x"00";
            when x"AFD" => q <= x"00";
            when x"AFE" => q <= x"00";
            when x"AFF" => q <= x"00";
            when x"B00" => q <= x"80";
            when x"B01" => q <= x"80";
            when x"B02" => q <= x"80";
            when x"B03" => q <= x"80";
            when x"B04" => q <= x"80";
            when x"B05" => q <= x"80";
            when x"B06" => q <= x"80";
            when x"B07" => q <= x"B8";
            when x"B08" => q <= x"B8";
            when x"B09" => q <= x"B8";
            when x"B0A" => q <= x"00";
            when x"B0B" => q <= x"00";
            when x"B0C" => q <= x"00";
            when x"B0D" => q <= x"00";
            when x"B0E" => q <= x"00";
            when x"B0F" => q <= x"00";
            when x"B10" => q <= x"B8";
            when x"B11" => q <= x"B8";
            when x"B12" => q <= x"B8";
            when x"B13" => q <= x"80";
            when x"B14" => q <= x"80";
            when x"B15" => q <= x"80";
            when x"B16" => q <= x"80";
            when x"B17" => q <= x"B8";
            when x"B18" => q <= x"B8";
            when x"B19" => q <= x"B8";
            when x"B1A" => q <= x"00";
            when x"B1B" => q <= x"00";
            when x"B1C" => q <= x"00";
            when x"B1D" => q <= x"00";
            when x"B1E" => q <= x"00";
            when x"B1F" => q <= x"00";
            when x"B20" => q <= x"87";
            when x"B21" => q <= x"87";
            when x"B22" => q <= x"87";
            when x"B23" => q <= x"80";
            when x"B24" => q <= x"80";
            when x"B25" => q <= x"80";
            when x"B26" => q <= x"80";
            when x"B27" => q <= x"B8";
            when x"B28" => q <= x"B8";
            when x"B29" => q <= x"B8";
            when x"B2A" => q <= x"00";
            when x"B2B" => q <= x"00";
            when x"B2C" => q <= x"00";
            when x"B2D" => q <= x"00";
            when x"B2E" => q <= x"00";
            when x"B2F" => q <= x"00";
            when x"B30" => q <= x"BF";
            when x"B31" => q <= x"BF";
            when x"B32" => q <= x"BF";
            when x"B33" => q <= x"80";
            when x"B34" => q <= x"80";
            when x"B35" => q <= x"80";
            when x"B36" => q <= x"80";
            when x"B37" => q <= x"B8";
            when x"B38" => q <= x"B8";
            when x"B39" => q <= x"B8";
            when x"B3A" => q <= x"00";
            when x"B3B" => q <= x"00";
            when x"B3C" => q <= x"00";
            when x"B3D" => q <= x"00";
            when x"B3E" => q <= x"00";
            when x"B3F" => q <= x"00";
            when x"B40" => q <= x"80";
            when x"B41" => q <= x"80";
            when x"B42" => q <= x"80";
            when x"B43" => q <= x"B8";
            when x"B44" => q <= x"B8";
            when x"B45" => q <= x"B8";
            when x"B46" => q <= x"B8";
            when x"B47" => q <= x"B8";
            when x"B48" => q <= x"B8";
            when x"B49" => q <= x"B8";
            when x"B4A" => q <= x"00";
            when x"B4B" => q <= x"00";
            when x"B4C" => q <= x"00";
            when x"B4D" => q <= x"00";
            when x"B4E" => q <= x"00";
            when x"B4F" => q <= x"00";
            when x"B50" => q <= x"B8";
            when x"B51" => q <= x"B8";
            when x"B52" => q <= x"B8";
            when x"B53" => q <= x"B8";
            when x"B54" => q <= x"B8";
            when x"B55" => q <= x"B8";
            when x"B56" => q <= x"B8";
            when x"B57" => q <= x"B8";
            when x"B58" => q <= x"B8";
            when x"B59" => q <= x"B8";
            when x"B5A" => q <= x"00";
            when x"B5B" => q <= x"00";
            when x"B5C" => q <= x"00";
            when x"B5D" => q <= x"00";
            when x"B5E" => q <= x"00";
            when x"B5F" => q <= x"00";
            when x"B60" => q <= x"87";
            when x"B61" => q <= x"87";
            when x"B62" => q <= x"87";
            when x"B63" => q <= x"B8";
            when x"B64" => q <= x"B8";
            when x"B65" => q <= x"B8";
            when x"B66" => q <= x"B8";
            when x"B67" => q <= x"B8";
            when x"B68" => q <= x"B8";
            when x"B69" => q <= x"B8";
            when x"B6A" => q <= x"00";
            when x"B6B" => q <= x"00";
            when x"B6C" => q <= x"00";
            when x"B6D" => q <= x"00";
            when x"B6E" => q <= x"00";
            when x"B6F" => q <= x"00";
            when x"B70" => q <= x"BF";
            when x"B71" => q <= x"BF";
            when x"B72" => q <= x"BF";
            when x"B73" => q <= x"B8";
            when x"B74" => q <= x"B8";
            when x"B75" => q <= x"B8";
            when x"B76" => q <= x"B8";
            when x"B77" => q <= x"B8";
            when x"B78" => q <= x"B8";
            when x"B79" => q <= x"B8";
            when x"B7A" => q <= x"00";
            when x"B7B" => q <= x"00";
            when x"B7C" => q <= x"00";
            when x"B7D" => q <= x"00";
            when x"B7E" => q <= x"00";
            when x"B7F" => q <= x"00";
            when x"B80" => q <= x"80";
            when x"B81" => q <= x"80";
            when x"B82" => q <= x"80";
            when x"B83" => q <= x"87";
            when x"B84" => q <= x"87";
            when x"B85" => q <= x"87";
            when x"B86" => q <= x"87";
            when x"B87" => q <= x"B8";
            when x"B88" => q <= x"B8";
            when x"B89" => q <= x"B8";
            when x"B8A" => q <= x"00";
            when x"B8B" => q <= x"00";
            when x"B8C" => q <= x"00";
            when x"B8D" => q <= x"00";
            when x"B8E" => q <= x"00";
            when x"B8F" => q <= x"00";
            when x"B90" => q <= x"B8";
            when x"B91" => q <= x"B8";
            when x"B92" => q <= x"B8";
            when x"B93" => q <= x"87";
            when x"B94" => q <= x"87";
            when x"B95" => q <= x"87";
            when x"B96" => q <= x"87";
            when x"B97" => q <= x"B8";
            when x"B98" => q <= x"B8";
            when x"B99" => q <= x"B8";
            when x"B9A" => q <= x"00";
            when x"B9B" => q <= x"00";
            when x"B9C" => q <= x"00";
            when x"B9D" => q <= x"00";
            when x"B9E" => q <= x"00";
            when x"B9F" => q <= x"00";
            when x"BA0" => q <= x"87";
            when x"BA1" => q <= x"87";
            when x"BA2" => q <= x"87";
            when x"BA3" => q <= x"87";
            when x"BA4" => q <= x"87";
            when x"BA5" => q <= x"87";
            when x"BA6" => q <= x"87";
            when x"BA7" => q <= x"B8";
            when x"BA8" => q <= x"B8";
            when x"BA9" => q <= x"B8";
            when x"BAA" => q <= x"00";
            when x"BAB" => q <= x"00";
            when x"BAC" => q <= x"00";
            when x"BAD" => q <= x"00";
            when x"BAE" => q <= x"00";
            when x"BAF" => q <= x"00";
            when x"BB0" => q <= x"BF";
            when x"BB1" => q <= x"BF";
            when x"BB2" => q <= x"BF";
            when x"BB3" => q <= x"87";
            when x"BB4" => q <= x"87";
            when x"BB5" => q <= x"87";
            when x"BB6" => q <= x"87";
            when x"BB7" => q <= x"B8";
            when x"BB8" => q <= x"B8";
            when x"BB9" => q <= x"B8";
            when x"BBA" => q <= x"00";
            when x"BBB" => q <= x"00";
            when x"BBC" => q <= x"00";
            when x"BBD" => q <= x"00";
            when x"BBE" => q <= x"00";
            when x"BBF" => q <= x"00";
            when x"BC0" => q <= x"80";
            when x"BC1" => q <= x"80";
            when x"BC2" => q <= x"80";
            when x"BC3" => q <= x"BF";
            when x"BC4" => q <= x"BF";
            when x"BC5" => q <= x"BF";
            when x"BC6" => q <= x"BF";
            when x"BC7" => q <= x"B8";
            when x"BC8" => q <= x"B8";
            when x"BC9" => q <= x"B8";
            when x"BCA" => q <= x"00";
            when x"BCB" => q <= x"00";
            when x"BCC" => q <= x"00";
            when x"BCD" => q <= x"00";
            when x"BCE" => q <= x"00";
            when x"BCF" => q <= x"00";
            when x"BD0" => q <= x"B8";
            when x"BD1" => q <= x"B8";
            when x"BD2" => q <= x"B8";
            when x"BD3" => q <= x"BF";
            when x"BD4" => q <= x"BF";
            when x"BD5" => q <= x"BF";
            when x"BD6" => q <= x"BF";
            when x"BD7" => q <= x"B8";
            when x"BD8" => q <= x"B8";
            when x"BD9" => q <= x"B8";
            when x"BDA" => q <= x"00";
            when x"BDB" => q <= x"00";
            when x"BDC" => q <= x"00";
            when x"BDD" => q <= x"00";
            when x"BDE" => q <= x"00";
            when x"BDF" => q <= x"00";
            when x"BE0" => q <= x"87";
            when x"BE1" => q <= x"87";
            when x"BE2" => q <= x"87";
            when x"BE3" => q <= x"BF";
            when x"BE4" => q <= x"BF";
            when x"BE5" => q <= x"BF";
            when x"BE6" => q <= x"BF";
            when x"BE7" => q <= x"B8";
            when x"BE8" => q <= x"B8";
            when x"BE9" => q <= x"B8";
            when x"BEA" => q <= x"00";
            when x"BEB" => q <= x"00";
            when x"BEC" => q <= x"00";
            when x"BED" => q <= x"00";
            when x"BEE" => q <= x"00";
            when x"BEF" => q <= x"00";
            when x"BF0" => q <= x"BF";
            when x"BF1" => q <= x"BF";
            when x"BF2" => q <= x"BF";
            when x"BF3" => q <= x"BF";
            when x"BF4" => q <= x"BF";
            when x"BF5" => q <= x"BF";
            when x"BF6" => q <= x"BF";
            when x"BF7" => q <= x"B8";
            when x"BF8" => q <= x"B8";
            when x"BF9" => q <= x"B8";
            when x"BFA" => q <= x"00";
            when x"BFB" => q <= x"00";
            when x"BFC" => q <= x"00";
            when x"BFD" => q <= x"00";
            when x"BFE" => q <= x"00";
            when x"BFF" => q <= x"00";
            when x"C00" => q <= x"00";
            when x"C01" => q <= x"0E";
            when x"C02" => q <= x"11";
            when x"C03" => q <= x"17";
            when x"C04" => q <= x"15";
            when x"C05" => q <= x"17";
            when x"C06" => q <= x"10";
            when x"C07" => q <= x"0E";
            when x"C08" => q <= x"00";
            when x"C09" => q <= x"00";
            when x"C0A" => q <= x"00";
            when x"C0B" => q <= x"00";
            when x"C0C" => q <= x"00";
            when x"C0D" => q <= x"00";
            when x"C0E" => q <= x"00";
            when x"C0F" => q <= x"00";
            when x"C10" => q <= x"00";
            when x"C11" => q <= x"04";
            when x"C12" => q <= x"0A";
            when x"C13" => q <= x"11";
            when x"C14" => q <= x"11";
            when x"C15" => q <= x"1F";
            when x"C16" => q <= x"11";
            when x"C17" => q <= x"11";
            when x"C18" => q <= x"00";
            when x"C19" => q <= x"00";
            when x"C1A" => q <= x"00";
            when x"C1B" => q <= x"00";
            when x"C1C" => q <= x"00";
            when x"C1D" => q <= x"00";
            when x"C1E" => q <= x"00";
            when x"C1F" => q <= x"00";
            when x"C20" => q <= x"00";
            when x"C21" => q <= x"1E";
            when x"C22" => q <= x"11";
            when x"C23" => q <= x"11";
            when x"C24" => q <= x"1E";
            when x"C25" => q <= x"11";
            when x"C26" => q <= x"11";
            when x"C27" => q <= x"1E";
            when x"C28" => q <= x"00";
            when x"C29" => q <= x"00";
            when x"C2A" => q <= x"00";
            when x"C2B" => q <= x"00";
            when x"C2C" => q <= x"00";
            when x"C2D" => q <= x"00";
            when x"C2E" => q <= x"00";
            when x"C2F" => q <= x"00";
            when x"C30" => q <= x"00";
            when x"C31" => q <= x"0E";
            when x"C32" => q <= x"11";
            when x"C33" => q <= x"10";
            when x"C34" => q <= x"10";
            when x"C35" => q <= x"10";
            when x"C36" => q <= x"11";
            when x"C37" => q <= x"0E";
            when x"C38" => q <= x"00";
            when x"C39" => q <= x"00";
            when x"C3A" => q <= x"00";
            when x"C3B" => q <= x"00";
            when x"C3C" => q <= x"00";
            when x"C3D" => q <= x"00";
            when x"C3E" => q <= x"00";
            when x"C3F" => q <= x"00";
            when x"C40" => q <= x"00";
            when x"C41" => q <= x"1E";
            when x"C42" => q <= x"11";
            when x"C43" => q <= x"11";
            when x"C44" => q <= x"11";
            when x"C45" => q <= x"11";
            when x"C46" => q <= x"11";
            when x"C47" => q <= x"1E";
            when x"C48" => q <= x"00";
            when x"C49" => q <= x"00";
            when x"C4A" => q <= x"00";
            when x"C4B" => q <= x"00";
            when x"C4C" => q <= x"00";
            when x"C4D" => q <= x"00";
            when x"C4E" => q <= x"00";
            when x"C4F" => q <= x"00";
            when x"C50" => q <= x"00";
            when x"C51" => q <= x"1F";
            when x"C52" => q <= x"10";
            when x"C53" => q <= x"10";
            when x"C54" => q <= x"1E";
            when x"C55" => q <= x"10";
            when x"C56" => q <= x"10";
            when x"C57" => q <= x"1F";
            when x"C58" => q <= x"00";
            when x"C59" => q <= x"00";
            when x"C5A" => q <= x"00";
            when x"C5B" => q <= x"00";
            when x"C5C" => q <= x"00";
            when x"C5D" => q <= x"00";
            when x"C5E" => q <= x"00";
            when x"C5F" => q <= x"00";
            when x"C60" => q <= x"00";
            when x"C61" => q <= x"1F";
            when x"C62" => q <= x"10";
            when x"C63" => q <= x"10";
            when x"C64" => q <= x"1E";
            when x"C65" => q <= x"10";
            when x"C66" => q <= x"10";
            when x"C67" => q <= x"10";
            when x"C68" => q <= x"00";
            when x"C69" => q <= x"00";
            when x"C6A" => q <= x"00";
            when x"C6B" => q <= x"00";
            when x"C6C" => q <= x"00";
            when x"C6D" => q <= x"00";
            when x"C6E" => q <= x"00";
            when x"C6F" => q <= x"00";
            when x"C70" => q <= x"00";
            when x"C71" => q <= x"0E";
            when x"C72" => q <= x"11";
            when x"C73" => q <= x"10";
            when x"C74" => q <= x"10";
            when x"C75" => q <= x"13";
            when x"C76" => q <= x"11";
            when x"C77" => q <= x"0F";
            when x"C78" => q <= x"00";
            when x"C79" => q <= x"00";
            when x"C7A" => q <= x"00";
            when x"C7B" => q <= x"00";
            when x"C7C" => q <= x"00";
            when x"C7D" => q <= x"00";
            when x"C7E" => q <= x"00";
            when x"C7F" => q <= x"00";
            when x"C80" => q <= x"00";
            when x"C81" => q <= x"11";
            when x"C82" => q <= x"11";
            when x"C83" => q <= x"11";
            when x"C84" => q <= x"1F";
            when x"C85" => q <= x"11";
            when x"C86" => q <= x"11";
            when x"C87" => q <= x"11";
            when x"C88" => q <= x"00";
            when x"C89" => q <= x"00";
            when x"C8A" => q <= x"00";
            when x"C8B" => q <= x"00";
            when x"C8C" => q <= x"00";
            when x"C8D" => q <= x"00";
            when x"C8E" => q <= x"00";
            when x"C8F" => q <= x"00";
            when x"C90" => q <= x"00";
            when x"C91" => q <= x"0E";
            when x"C92" => q <= x"04";
            when x"C93" => q <= x"04";
            when x"C94" => q <= x"04";
            when x"C95" => q <= x"04";
            when x"C96" => q <= x"04";
            when x"C97" => q <= x"0E";
            when x"C98" => q <= x"00";
            when x"C99" => q <= x"00";
            when x"C9A" => q <= x"00";
            when x"C9B" => q <= x"00";
            when x"C9C" => q <= x"00";
            when x"C9D" => q <= x"00";
            when x"C9E" => q <= x"00";
            when x"C9F" => q <= x"00";
            when x"CA0" => q <= x"00";
            when x"CA1" => q <= x"01";
            when x"CA2" => q <= x"01";
            when x"CA3" => q <= x"01";
            when x"CA4" => q <= x"01";
            when x"CA5" => q <= x"01";
            when x"CA6" => q <= x"11";
            when x"CA7" => q <= x"0E";
            when x"CA8" => q <= x"00";
            when x"CA9" => q <= x"00";
            when x"CAA" => q <= x"00";
            when x"CAB" => q <= x"00";
            when x"CAC" => q <= x"00";
            when x"CAD" => q <= x"00";
            when x"CAE" => q <= x"00";
            when x"CAF" => q <= x"00";
            when x"CB0" => q <= x"00";
            when x"CB1" => q <= x"11";
            when x"CB2" => q <= x"12";
            when x"CB3" => q <= x"14";
            when x"CB4" => q <= x"18";
            when x"CB5" => q <= x"14";
            when x"CB6" => q <= x"12";
            when x"CB7" => q <= x"11";
            when x"CB8" => q <= x"00";
            when x"CB9" => q <= x"00";
            when x"CBA" => q <= x"00";
            when x"CBB" => q <= x"00";
            when x"CBC" => q <= x"00";
            when x"CBD" => q <= x"00";
            when x"CBE" => q <= x"00";
            when x"CBF" => q <= x"00";
            when x"CC0" => q <= x"00";
            when x"CC1" => q <= x"10";
            when x"CC2" => q <= x"10";
            when x"CC3" => q <= x"10";
            when x"CC4" => q <= x"10";
            when x"CC5" => q <= x"10";
            when x"CC6" => q <= x"10";
            when x"CC7" => q <= x"1F";
            when x"CC8" => q <= x"00";
            when x"CC9" => q <= x"00";
            when x"CCA" => q <= x"00";
            when x"CCB" => q <= x"00";
            when x"CCC" => q <= x"00";
            when x"CCD" => q <= x"00";
            when x"CCE" => q <= x"00";
            when x"CCF" => q <= x"00";
            when x"CD0" => q <= x"00";
            when x"CD1" => q <= x"11";
            when x"CD2" => q <= x"1B";
            when x"CD3" => q <= x"15";
            when x"CD4" => q <= x"15";
            when x"CD5" => q <= x"11";
            when x"CD6" => q <= x"11";
            when x"CD7" => q <= x"11";
            when x"CD8" => q <= x"00";
            when x"CD9" => q <= x"00";
            when x"CDA" => q <= x"00";
            when x"CDB" => q <= x"00";
            when x"CDC" => q <= x"00";
            when x"CDD" => q <= x"00";
            when x"CDE" => q <= x"00";
            when x"CDF" => q <= x"00";
            when x"CE0" => q <= x"00";
            when x"CE1" => q <= x"11";
            when x"CE2" => q <= x"11";
            when x"CE3" => q <= x"19";
            when x"CE4" => q <= x"15";
            when x"CE5" => q <= x"13";
            when x"CE6" => q <= x"11";
            when x"CE7" => q <= x"11";
            when x"CE8" => q <= x"00";
            when x"CE9" => q <= x"00";
            when x"CEA" => q <= x"00";
            when x"CEB" => q <= x"00";
            when x"CEC" => q <= x"00";
            when x"CED" => q <= x"00";
            when x"CEE" => q <= x"00";
            when x"CEF" => q <= x"00";
            when x"CF0" => q <= x"00";
            when x"CF1" => q <= x"0E";
            when x"CF2" => q <= x"11";
            when x"CF3" => q <= x"11";
            when x"CF4" => q <= x"11";
            when x"CF5" => q <= x"11";
            when x"CF6" => q <= x"11";
            when x"CF7" => q <= x"0E";
            when x"CF8" => q <= x"00";
            when x"CF9" => q <= x"00";
            when x"CFA" => q <= x"00";
            when x"CFB" => q <= x"00";
            when x"CFC" => q <= x"00";
            when x"CFD" => q <= x"00";
            when x"CFE" => q <= x"00";
            when x"CFF" => q <= x"00";
            when x"D00" => q <= x"00";
            when x"D01" => q <= x"1E";
            when x"D02" => q <= x"11";
            when x"D03" => q <= x"11";
            when x"D04" => q <= x"1E";
            when x"D05" => q <= x"10";
            when x"D06" => q <= x"10";
            when x"D07" => q <= x"10";
            when x"D08" => q <= x"00";
            when x"D09" => q <= x"00";
            when x"D0A" => q <= x"00";
            when x"D0B" => q <= x"00";
            when x"D0C" => q <= x"00";
            when x"D0D" => q <= x"00";
            when x"D0E" => q <= x"00";
            when x"D0F" => q <= x"00";
            when x"D10" => q <= x"00";
            when x"D11" => q <= x"0E";
            when x"D12" => q <= x"11";
            when x"D13" => q <= x"11";
            when x"D14" => q <= x"11";
            when x"D15" => q <= x"15";
            when x"D16" => q <= x"12";
            when x"D17" => q <= x"0D";
            when x"D18" => q <= x"00";
            when x"D19" => q <= x"00";
            when x"D1A" => q <= x"00";
            when x"D1B" => q <= x"00";
            when x"D1C" => q <= x"00";
            when x"D1D" => q <= x"00";
            when x"D1E" => q <= x"00";
            when x"D1F" => q <= x"00";
            when x"D20" => q <= x"00";
            when x"D21" => q <= x"1E";
            when x"D22" => q <= x"11";
            when x"D23" => q <= x"11";
            when x"D24" => q <= x"1E";
            when x"D25" => q <= x"14";
            when x"D26" => q <= x"12";
            when x"D27" => q <= x"11";
            when x"D28" => q <= x"00";
            when x"D29" => q <= x"00";
            when x"D2A" => q <= x"00";
            when x"D2B" => q <= x"00";
            when x"D2C" => q <= x"00";
            when x"D2D" => q <= x"00";
            when x"D2E" => q <= x"00";
            when x"D2F" => q <= x"00";
            when x"D30" => q <= x"00";
            when x"D31" => q <= x"0E";
            when x"D32" => q <= x"11";
            when x"D33" => q <= x"10";
            when x"D34" => q <= x"0E";
            when x"D35" => q <= x"01";
            when x"D36" => q <= x"11";
            when x"D37" => q <= x"0E";
            when x"D38" => q <= x"00";
            when x"D39" => q <= x"00";
            when x"D3A" => q <= x"00";
            when x"D3B" => q <= x"00";
            when x"D3C" => q <= x"00";
            when x"D3D" => q <= x"00";
            when x"D3E" => q <= x"00";
            when x"D3F" => q <= x"00";
            when x"D40" => q <= x"00";
            when x"D41" => q <= x"1F";
            when x"D42" => q <= x"04";
            when x"D43" => q <= x"04";
            when x"D44" => q <= x"04";
            when x"D45" => q <= x"04";
            when x"D46" => q <= x"04";
            when x"D47" => q <= x"04";
            when x"D48" => q <= x"00";
            when x"D49" => q <= x"00";
            when x"D4A" => q <= x"00";
            when x"D4B" => q <= x"00";
            when x"D4C" => q <= x"00";
            when x"D4D" => q <= x"00";
            when x"D4E" => q <= x"00";
            when x"D4F" => q <= x"00";
            when x"D50" => q <= x"00";
            when x"D51" => q <= x"11";
            when x"D52" => q <= x"11";
            when x"D53" => q <= x"11";
            when x"D54" => q <= x"11";
            when x"D55" => q <= x"11";
            when x"D56" => q <= x"11";
            when x"D57" => q <= x"0E";
            when x"D58" => q <= x"00";
            when x"D59" => q <= x"00";
            when x"D5A" => q <= x"00";
            when x"D5B" => q <= x"00";
            when x"D5C" => q <= x"00";
            when x"D5D" => q <= x"00";
            when x"D5E" => q <= x"00";
            when x"D5F" => q <= x"00";
            when x"D60" => q <= x"00";
            when x"D61" => q <= x"11";
            when x"D62" => q <= x"11";
            when x"D63" => q <= x"11";
            when x"D64" => q <= x"0A";
            when x"D65" => q <= x"0A";
            when x"D66" => q <= x"04";
            when x"D67" => q <= x"04";
            when x"D68" => q <= x"00";
            when x"D69" => q <= x"00";
            when x"D6A" => q <= x"00";
            when x"D6B" => q <= x"00";
            when x"D6C" => q <= x"00";
            when x"D6D" => q <= x"00";
            when x"D6E" => q <= x"00";
            when x"D6F" => q <= x"00";
            when x"D70" => q <= x"00";
            when x"D71" => q <= x"11";
            when x"D72" => q <= x"11";
            when x"D73" => q <= x"11";
            when x"D74" => q <= x"15";
            when x"D75" => q <= x"15";
            when x"D76" => q <= x"15";
            when x"D77" => q <= x"0A";
            when x"D78" => q <= x"00";
            when x"D79" => q <= x"00";
            when x"D7A" => q <= x"00";
            when x"D7B" => q <= x"00";
            when x"D7C" => q <= x"00";
            when x"D7D" => q <= x"00";
            when x"D7E" => q <= x"00";
            when x"D7F" => q <= x"00";
            when x"D80" => q <= x"00";
            when x"D81" => q <= x"11";
            when x"D82" => q <= x"11";
            when x"D83" => q <= x"0A";
            when x"D84" => q <= x"04";
            when x"D85" => q <= x"0A";
            when x"D86" => q <= x"11";
            when x"D87" => q <= x"11";
            when x"D88" => q <= x"00";
            when x"D89" => q <= x"00";
            when x"D8A" => q <= x"00";
            when x"D8B" => q <= x"00";
            when x"D8C" => q <= x"00";
            when x"D8D" => q <= x"00";
            when x"D8E" => q <= x"00";
            when x"D8F" => q <= x"00";
            when x"D90" => q <= x"00";
            when x"D91" => q <= x"11";
            when x"D92" => q <= x"11";
            when x"D93" => q <= x"0A";
            when x"D94" => q <= x"04";
            when x"D95" => q <= x"04";
            when x"D96" => q <= x"04";
            when x"D97" => q <= x"04";
            when x"D98" => q <= x"00";
            when x"D99" => q <= x"00";
            when x"D9A" => q <= x"00";
            when x"D9B" => q <= x"00";
            when x"D9C" => q <= x"00";
            when x"D9D" => q <= x"00";
            when x"D9E" => q <= x"00";
            when x"D9F" => q <= x"00";
            when x"DA0" => q <= x"00";
            when x"DA1" => q <= x"1F";
            when x"DA2" => q <= x"01";
            when x"DA3" => q <= x"02";
            when x"DA4" => q <= x"04";
            when x"DA5" => q <= x"08";
            when x"DA6" => q <= x"10";
            when x"DA7" => q <= x"1F";
            when x"DA8" => q <= x"00";
            when x"DA9" => q <= x"00";
            when x"DAA" => q <= x"00";
            when x"DAB" => q <= x"00";
            when x"DAC" => q <= x"00";
            when x"DAD" => q <= x"00";
            when x"DAE" => q <= x"00";
            when x"DAF" => q <= x"00";
            when x"DB0" => q <= x"00";
            when x"DB1" => q <= x"00";
            when x"DB2" => q <= x"04";
            when x"DB3" => q <= x"08";
            when x"DB4" => q <= x"1F";
            when x"DB5" => q <= x"08";
            when x"DB6" => q <= x"04";
            when x"DB7" => q <= x"00";
            when x"DB8" => q <= x"00";
            when x"DB9" => q <= x"00";
            when x"DBA" => q <= x"00";
            when x"DBB" => q <= x"00";
            when x"DBC" => q <= x"00";
            when x"DBD" => q <= x"00";
            when x"DBE" => q <= x"00";
            when x"DBF" => q <= x"00";
            when x"DC0" => q <= x"00";
            when x"DC1" => q <= x"10";
            when x"DC2" => q <= x"10";
            when x"DC3" => q <= x"10";
            when x"DC4" => q <= x"10";
            when x"DC5" => q <= x"16";
            when x"DC6" => q <= x"01";
            when x"DC7" => q <= x"02";
            when x"DC8" => q <= x"04";
            when x"DC9" => q <= x"07";
            when x"DCA" => q <= x"00";
            when x"DCB" => q <= x"00";
            when x"DCC" => q <= x"00";
            when x"DCD" => q <= x"00";
            when x"DCE" => q <= x"00";
            when x"DCF" => q <= x"00";
            when x"DD0" => q <= x"00";
            when x"DD1" => q <= x"00";
            when x"DD2" => q <= x"04";
            when x"DD3" => q <= x"02";
            when x"DD4" => q <= x"1F";
            when x"DD5" => q <= x"02";
            when x"DD6" => q <= x"04";
            when x"DD7" => q <= x"00";
            when x"DD8" => q <= x"00";
            when x"DD9" => q <= x"00";
            when x"DDA" => q <= x"00";
            when x"DDB" => q <= x"00";
            when x"DDC" => q <= x"00";
            when x"DDD" => q <= x"00";
            when x"DDE" => q <= x"00";
            when x"DDF" => q <= x"00";
            when x"DE0" => q <= x"00";
            when x"DE1" => q <= x"00";
            when x"DE2" => q <= x"04";
            when x"DE3" => q <= x"0E";
            when x"DE4" => q <= x"15";
            when x"DE5" => q <= x"04";
            when x"DE6" => q <= x"04";
            when x"DE7" => q <= x"00";
            when x"DE8" => q <= x"00";
            when x"DE9" => q <= x"00";
            when x"DEA" => q <= x"00";
            when x"DEB" => q <= x"00";
            when x"DEC" => q <= x"00";
            when x"DED" => q <= x"00";
            when x"DEE" => q <= x"00";
            when x"DEF" => q <= x"00";
            when x"DF0" => q <= x"00";
            when x"DF1" => q <= x"0A";
            when x"DF2" => q <= x"0A";
            when x"DF3" => q <= x"1F";
            when x"DF4" => q <= x"0A";
            when x"DF5" => q <= x"1F";
            when x"DF6" => q <= x"0A";
            when x"DF7" => q <= x"0A";
            when x"DF8" => q <= x"00";
            when x"DF9" => q <= x"00";
            when x"DFA" => q <= x"00";
            when x"DFB" => q <= x"00";
            when x"DFC" => q <= x"00";
            when x"DFD" => q <= x"00";
            when x"DFE" => q <= x"00";
            when x"DFF" => q <= x"00";
            when x"E00" => q <= x"80";
            when x"E01" => q <= x"80";
            when x"E02" => q <= x"80";
            when x"E03" => q <= x"80";
            when x"E04" => q <= x"80";
            when x"E05" => q <= x"80";
            when x"E06" => q <= x"80";
            when x"E07" => q <= x"87";
            when x"E08" => q <= x"87";
            when x"E09" => q <= x"87";
            when x"E0A" => q <= x"00";
            when x"E0B" => q <= x"00";
            when x"E0C" => q <= x"00";
            when x"E0D" => q <= x"00";
            when x"E0E" => q <= x"00";
            when x"E0F" => q <= x"00";
            when x"E10" => q <= x"B8";
            when x"E11" => q <= x"B8";
            when x"E12" => q <= x"B8";
            when x"E13" => q <= x"80";
            when x"E14" => q <= x"80";
            when x"E15" => q <= x"80";
            when x"E16" => q <= x"80";
            when x"E17" => q <= x"87";
            when x"E18" => q <= x"87";
            when x"E19" => q <= x"87";
            when x"E1A" => q <= x"00";
            when x"E1B" => q <= x"00";
            when x"E1C" => q <= x"00";
            when x"E1D" => q <= x"00";
            when x"E1E" => q <= x"00";
            when x"E1F" => q <= x"00";
            when x"E20" => q <= x"87";
            when x"E21" => q <= x"87";
            when x"E22" => q <= x"87";
            when x"E23" => q <= x"80";
            when x"E24" => q <= x"80";
            when x"E25" => q <= x"80";
            when x"E26" => q <= x"80";
            when x"E27" => q <= x"87";
            when x"E28" => q <= x"87";
            when x"E29" => q <= x"87";
            when x"E2A" => q <= x"00";
            when x"E2B" => q <= x"00";
            when x"E2C" => q <= x"00";
            when x"E2D" => q <= x"00";
            when x"E2E" => q <= x"00";
            when x"E2F" => q <= x"00";
            when x"E30" => q <= x"BF";
            when x"E31" => q <= x"BF";
            when x"E32" => q <= x"BF";
            when x"E33" => q <= x"80";
            when x"E34" => q <= x"80";
            when x"E35" => q <= x"80";
            when x"E36" => q <= x"80";
            when x"E37" => q <= x"87";
            when x"E38" => q <= x"87";
            when x"E39" => q <= x"87";
            when x"E3A" => q <= x"00";
            when x"E3B" => q <= x"00";
            when x"E3C" => q <= x"00";
            when x"E3D" => q <= x"00";
            when x"E3E" => q <= x"00";
            when x"E3F" => q <= x"00";
            when x"E40" => q <= x"80";
            when x"E41" => q <= x"80";
            when x"E42" => q <= x"80";
            when x"E43" => q <= x"B8";
            when x"E44" => q <= x"B8";
            when x"E45" => q <= x"B8";
            when x"E46" => q <= x"B8";
            when x"E47" => q <= x"87";
            when x"E48" => q <= x"87";
            when x"E49" => q <= x"87";
            when x"E4A" => q <= x"00";
            when x"E4B" => q <= x"00";
            when x"E4C" => q <= x"00";
            when x"E4D" => q <= x"00";
            when x"E4E" => q <= x"00";
            when x"E4F" => q <= x"00";
            when x"E50" => q <= x"B8";
            when x"E51" => q <= x"B8";
            when x"E52" => q <= x"B8";
            when x"E53" => q <= x"B8";
            when x"E54" => q <= x"B8";
            when x"E55" => q <= x"B8";
            when x"E56" => q <= x"B8";
            when x"E57" => q <= x"87";
            when x"E58" => q <= x"87";
            when x"E59" => q <= x"87";
            when x"E5A" => q <= x"00";
            when x"E5B" => q <= x"00";
            when x"E5C" => q <= x"00";
            when x"E5D" => q <= x"00";
            when x"E5E" => q <= x"00";
            when x"E5F" => q <= x"00";
            when x"E60" => q <= x"87";
            when x"E61" => q <= x"87";
            when x"E62" => q <= x"87";
            when x"E63" => q <= x"B8";
            when x"E64" => q <= x"B8";
            when x"E65" => q <= x"B8";
            when x"E66" => q <= x"B8";
            when x"E67" => q <= x"87";
            when x"E68" => q <= x"87";
            when x"E69" => q <= x"87";
            when x"E6A" => q <= x"00";
            when x"E6B" => q <= x"00";
            when x"E6C" => q <= x"00";
            when x"E6D" => q <= x"00";
            when x"E6E" => q <= x"00";
            when x"E6F" => q <= x"00";
            when x"E70" => q <= x"BF";
            when x"E71" => q <= x"BF";
            when x"E72" => q <= x"BF";
            when x"E73" => q <= x"B8";
            when x"E74" => q <= x"B8";
            when x"E75" => q <= x"B8";
            when x"E76" => q <= x"B8";
            when x"E77" => q <= x"87";
            when x"E78" => q <= x"87";
            when x"E79" => q <= x"87";
            when x"E7A" => q <= x"00";
            when x"E7B" => q <= x"00";
            when x"E7C" => q <= x"00";
            when x"E7D" => q <= x"00";
            when x"E7E" => q <= x"00";
            when x"E7F" => q <= x"00";
            when x"E80" => q <= x"80";
            when x"E81" => q <= x"80";
            when x"E82" => q <= x"80";
            when x"E83" => q <= x"87";
            when x"E84" => q <= x"87";
            when x"E85" => q <= x"87";
            when x"E86" => q <= x"87";
            when x"E87" => q <= x"87";
            when x"E88" => q <= x"87";
            when x"E89" => q <= x"87";
            when x"E8A" => q <= x"00";
            when x"E8B" => q <= x"00";
            when x"E8C" => q <= x"00";
            when x"E8D" => q <= x"00";
            when x"E8E" => q <= x"00";
            when x"E8F" => q <= x"00";
            when x"E90" => q <= x"B8";
            when x"E91" => q <= x"B8";
            when x"E92" => q <= x"B8";
            when x"E93" => q <= x"87";
            when x"E94" => q <= x"87";
            when x"E95" => q <= x"87";
            when x"E96" => q <= x"87";
            when x"E97" => q <= x"87";
            when x"E98" => q <= x"87";
            when x"E99" => q <= x"87";
            when x"E9A" => q <= x"00";
            when x"E9B" => q <= x"00";
            when x"E9C" => q <= x"00";
            when x"E9D" => q <= x"00";
            when x"E9E" => q <= x"00";
            when x"E9F" => q <= x"00";
            when x"EA0" => q <= x"87";
            when x"EA1" => q <= x"87";
            when x"EA2" => q <= x"87";
            when x"EA3" => q <= x"87";
            when x"EA4" => q <= x"87";
            when x"EA5" => q <= x"87";
            when x"EA6" => q <= x"87";
            when x"EA7" => q <= x"87";
            when x"EA8" => q <= x"87";
            when x"EA9" => q <= x"87";
            when x"EAA" => q <= x"00";
            when x"EAB" => q <= x"00";
            when x"EAC" => q <= x"00";
            when x"EAD" => q <= x"00";
            when x"EAE" => q <= x"00";
            when x"EAF" => q <= x"00";
            when x"EB0" => q <= x"BF";
            when x"EB1" => q <= x"BF";
            when x"EB2" => q <= x"BF";
            when x"EB3" => q <= x"87";
            when x"EB4" => q <= x"87";
            when x"EB5" => q <= x"87";
            when x"EB6" => q <= x"87";
            when x"EB7" => q <= x"87";
            when x"EB8" => q <= x"87";
            when x"EB9" => q <= x"87";
            when x"EBA" => q <= x"00";
            when x"EBB" => q <= x"00";
            when x"EBC" => q <= x"00";
            when x"EBD" => q <= x"00";
            when x"EBE" => q <= x"00";
            when x"EBF" => q <= x"00";
            when x"EC0" => q <= x"80";
            when x"EC1" => q <= x"80";
            when x"EC2" => q <= x"80";
            when x"EC3" => q <= x"BF";
            when x"EC4" => q <= x"BF";
            when x"EC5" => q <= x"BF";
            when x"EC6" => q <= x"BF";
            when x"EC7" => q <= x"87";
            when x"EC8" => q <= x"87";
            when x"EC9" => q <= x"87";
            when x"ECA" => q <= x"00";
            when x"ECB" => q <= x"00";
            when x"ECC" => q <= x"00";
            when x"ECD" => q <= x"00";
            when x"ECE" => q <= x"00";
            when x"ECF" => q <= x"00";
            when x"ED0" => q <= x"B8";
            when x"ED1" => q <= x"B8";
            when x"ED2" => q <= x"B8";
            when x"ED3" => q <= x"BF";
            when x"ED4" => q <= x"BF";
            when x"ED5" => q <= x"BF";
            when x"ED6" => q <= x"BF";
            when x"ED7" => q <= x"87";
            when x"ED8" => q <= x"87";
            when x"ED9" => q <= x"87";
            when x"EDA" => q <= x"00";
            when x"EDB" => q <= x"00";
            when x"EDC" => q <= x"00";
            when x"EDD" => q <= x"00";
            when x"EDE" => q <= x"00";
            when x"EDF" => q <= x"00";
            when x"EE0" => q <= x"87";
            when x"EE1" => q <= x"87";
            when x"EE2" => q <= x"87";
            when x"EE3" => q <= x"BF";
            when x"EE4" => q <= x"BF";
            when x"EE5" => q <= x"BF";
            when x"EE6" => q <= x"BF";
            when x"EE7" => q <= x"87";
            when x"EE8" => q <= x"87";
            when x"EE9" => q <= x"87";
            when x"EEA" => q <= x"00";
            when x"EEB" => q <= x"00";
            when x"EEC" => q <= x"00";
            when x"EED" => q <= x"00";
            when x"EEE" => q <= x"00";
            when x"EEF" => q <= x"00";
            when x"EF0" => q <= x"BF";
            when x"EF1" => q <= x"BF";
            when x"EF2" => q <= x"BF";
            when x"EF3" => q <= x"BF";
            when x"EF4" => q <= x"BF";
            when x"EF5" => q <= x"BF";
            when x"EF6" => q <= x"BF";
            when x"EF7" => q <= x"87";
            when x"EF8" => q <= x"87";
            when x"EF9" => q <= x"87";
            when x"EFA" => q <= x"00";
            when x"EFB" => q <= x"00";
            when x"EFC" => q <= x"00";
            when x"EFD" => q <= x"00";
            when x"EFE" => q <= x"00";
            when x"EFF" => q <= x"00";
            when x"F00" => q <= x"80";
            when x"F01" => q <= x"80";
            when x"F02" => q <= x"80";
            when x"F03" => q <= x"80";
            when x"F04" => q <= x"80";
            when x"F05" => q <= x"80";
            when x"F06" => q <= x"80";
            when x"F07" => q <= x"BF";
            when x"F08" => q <= x"BF";
            when x"F09" => q <= x"BF";
            when x"F0A" => q <= x"00";
            when x"F0B" => q <= x"00";
            when x"F0C" => q <= x"00";
            when x"F0D" => q <= x"00";
            when x"F0E" => q <= x"00";
            when x"F0F" => q <= x"00";
            when x"F10" => q <= x"B8";
            when x"F11" => q <= x"B8";
            when x"F12" => q <= x"B8";
            when x"F13" => q <= x"80";
            when x"F14" => q <= x"80";
            when x"F15" => q <= x"80";
            when x"F16" => q <= x"80";
            when x"F17" => q <= x"BF";
            when x"F18" => q <= x"BF";
            when x"F19" => q <= x"BF";
            when x"F1A" => q <= x"00";
            when x"F1B" => q <= x"00";
            when x"F1C" => q <= x"00";
            when x"F1D" => q <= x"00";
            when x"F1E" => q <= x"00";
            when x"F1F" => q <= x"00";
            when x"F20" => q <= x"87";
            when x"F21" => q <= x"87";
            when x"F22" => q <= x"87";
            when x"F23" => q <= x"80";
            when x"F24" => q <= x"80";
            when x"F25" => q <= x"80";
            when x"F26" => q <= x"80";
            when x"F27" => q <= x"BF";
            when x"F28" => q <= x"BF";
            when x"F29" => q <= x"BF";
            when x"F2A" => q <= x"00";
            when x"F2B" => q <= x"00";
            when x"F2C" => q <= x"00";
            when x"F2D" => q <= x"00";
            when x"F2E" => q <= x"00";
            when x"F2F" => q <= x"00";
            when x"F30" => q <= x"BF";
            when x"F31" => q <= x"BF";
            when x"F32" => q <= x"BF";
            when x"F33" => q <= x"80";
            when x"F34" => q <= x"80";
            when x"F35" => q <= x"80";
            when x"F36" => q <= x"80";
            when x"F37" => q <= x"BF";
            when x"F38" => q <= x"BF";
            when x"F39" => q <= x"BF";
            when x"F3A" => q <= x"00";
            when x"F3B" => q <= x"00";
            when x"F3C" => q <= x"00";
            when x"F3D" => q <= x"00";
            when x"F3E" => q <= x"00";
            when x"F3F" => q <= x"00";
            when x"F40" => q <= x"80";
            when x"F41" => q <= x"80";
            when x"F42" => q <= x"80";
            when x"F43" => q <= x"B8";
            when x"F44" => q <= x"B8";
            when x"F45" => q <= x"B8";
            when x"F46" => q <= x"B8";
            when x"F47" => q <= x"BF";
            when x"F48" => q <= x"BF";
            when x"F49" => q <= x"BF";
            when x"F4A" => q <= x"00";
            when x"F4B" => q <= x"00";
            when x"F4C" => q <= x"00";
            when x"F4D" => q <= x"00";
            when x"F4E" => q <= x"00";
            when x"F4F" => q <= x"00";
            when x"F50" => q <= x"B8";
            when x"F51" => q <= x"B8";
            when x"F52" => q <= x"B8";
            when x"F53" => q <= x"B8";
            when x"F54" => q <= x"B8";
            when x"F55" => q <= x"B8";
            when x"F56" => q <= x"B8";
            when x"F57" => q <= x"BF";
            when x"F58" => q <= x"BF";
            when x"F59" => q <= x"BF";
            when x"F5A" => q <= x"00";
            when x"F5B" => q <= x"00";
            when x"F5C" => q <= x"00";
            when x"F5D" => q <= x"00";
            when x"F5E" => q <= x"00";
            when x"F5F" => q <= x"00";
            when x"F60" => q <= x"87";
            when x"F61" => q <= x"87";
            when x"F62" => q <= x"87";
            when x"F63" => q <= x"B8";
            when x"F64" => q <= x"B8";
            when x"F65" => q <= x"B8";
            when x"F66" => q <= x"B8";
            when x"F67" => q <= x"BF";
            when x"F68" => q <= x"BF";
            when x"F69" => q <= x"BF";
            when x"F6A" => q <= x"00";
            when x"F6B" => q <= x"00";
            when x"F6C" => q <= x"00";
            when x"F6D" => q <= x"00";
            when x"F6E" => q <= x"00";
            when x"F6F" => q <= x"00";
            when x"F70" => q <= x"BF";
            when x"F71" => q <= x"BF";
            when x"F72" => q <= x"BF";
            when x"F73" => q <= x"B8";
            when x"F74" => q <= x"B8";
            when x"F75" => q <= x"B8";
            when x"F76" => q <= x"B8";
            when x"F77" => q <= x"BF";
            when x"F78" => q <= x"BF";
            when x"F79" => q <= x"BF";
            when x"F7A" => q <= x"00";
            when x"F7B" => q <= x"00";
            when x"F7C" => q <= x"00";
            when x"F7D" => q <= x"00";
            when x"F7E" => q <= x"00";
            when x"F7F" => q <= x"00";
            when x"F80" => q <= x"80";
            when x"F81" => q <= x"80";
            when x"F82" => q <= x"80";
            when x"F83" => q <= x"87";
            when x"F84" => q <= x"87";
            when x"F85" => q <= x"87";
            when x"F86" => q <= x"87";
            when x"F87" => q <= x"BF";
            when x"F88" => q <= x"BF";
            when x"F89" => q <= x"BF";
            when x"F8A" => q <= x"00";
            when x"F8B" => q <= x"00";
            when x"F8C" => q <= x"00";
            when x"F8D" => q <= x"00";
            when x"F8E" => q <= x"00";
            when x"F8F" => q <= x"00";
            when x"F90" => q <= x"B8";
            when x"F91" => q <= x"B8";
            when x"F92" => q <= x"B8";
            when x"F93" => q <= x"87";
            when x"F94" => q <= x"87";
            when x"F95" => q <= x"87";
            when x"F96" => q <= x"87";
            when x"F97" => q <= x"BF";
            when x"F98" => q <= x"BF";
            when x"F99" => q <= x"BF";
            when x"F9A" => q <= x"00";
            when x"F9B" => q <= x"00";
            when x"F9C" => q <= x"00";
            when x"F9D" => q <= x"00";
            when x"F9E" => q <= x"00";
            when x"F9F" => q <= x"00";
            when x"FA0" => q <= x"87";
            when x"FA1" => q <= x"87";
            when x"FA2" => q <= x"87";
            when x"FA3" => q <= x"87";
            when x"FA4" => q <= x"87";
            when x"FA5" => q <= x"87";
            when x"FA6" => q <= x"87";
            when x"FA7" => q <= x"BF";
            when x"FA8" => q <= x"BF";
            when x"FA9" => q <= x"BF";
            when x"FAA" => q <= x"00";
            when x"FAB" => q <= x"00";
            when x"FAC" => q <= x"00";
            when x"FAD" => q <= x"00";
            when x"FAE" => q <= x"00";
            when x"FAF" => q <= x"00";
            when x"FB0" => q <= x"BF";
            when x"FB1" => q <= x"BF";
            when x"FB2" => q <= x"BF";
            when x"FB3" => q <= x"87";
            when x"FB4" => q <= x"87";
            when x"FB5" => q <= x"87";
            when x"FB6" => q <= x"87";
            when x"FB7" => q <= x"BF";
            when x"FB8" => q <= x"BF";
            when x"FB9" => q <= x"BF";
            when x"FBA" => q <= x"00";
            when x"FBB" => q <= x"00";
            when x"FBC" => q <= x"00";
            when x"FBD" => q <= x"00";
            when x"FBE" => q <= x"00";
            when x"FBF" => q <= x"00";
            when x"FC0" => q <= x"80";
            when x"FC1" => q <= x"80";
            when x"FC2" => q <= x"80";
            when x"FC3" => q <= x"BF";
            when x"FC4" => q <= x"BF";
            when x"FC5" => q <= x"BF";
            when x"FC6" => q <= x"BF";
            when x"FC7" => q <= x"BF";
            when x"FC8" => q <= x"BF";
            when x"FC9" => q <= x"BF";
            when x"FCA" => q <= x"00";
            when x"FCB" => q <= x"00";
            when x"FCC" => q <= x"00";
            when x"FCD" => q <= x"00";
            when x"FCE" => q <= x"00";
            when x"FCF" => q <= x"00";
            when x"FD0" => q <= x"B8";
            when x"FD1" => q <= x"B8";
            when x"FD2" => q <= x"B8";
            when x"FD3" => q <= x"BF";
            when x"FD4" => q <= x"BF";
            when x"FD5" => q <= x"BF";
            when x"FD6" => q <= x"BF";
            when x"FD7" => q <= x"BF";
            when x"FD8" => q <= x"BF";
            when x"FD9" => q <= x"BF";
            when x"FDA" => q <= x"00";
            when x"FDB" => q <= x"00";
            when x"FDC" => q <= x"00";
            when x"FDD" => q <= x"00";
            when x"FDE" => q <= x"00";
            when x"FDF" => q <= x"00";
            when x"FE0" => q <= x"87";
            when x"FE1" => q <= x"87";
            when x"FE2" => q <= x"87";
            when x"FE3" => q <= x"BF";
            when x"FE4" => q <= x"BF";
            when x"FE5" => q <= x"BF";
            when x"FE6" => q <= x"BF";
            when x"FE7" => q <= x"BF";
            when x"FE8" => q <= x"BF";
            when x"FE9" => q <= x"BF";
            when x"FEA" => q <= x"00";
            when x"FEB" => q <= x"00";
            when x"FEC" => q <= x"00";
            when x"FED" => q <= x"00";
            when x"FEE" => q <= x"00";
            when x"FEF" => q <= x"00";
            when x"FF0" => q <= x"BF";
            when x"FF1" => q <= x"BF";
            when x"FF2" => q <= x"BF";
            when x"FF3" => q <= x"BF";
            when x"FF4" => q <= x"BF";
            when x"FF5" => q <= x"BF";
            when x"FF6" => q <= x"BF";
            when x"FF7" => q <= x"BF";
            when x"FF8" => q <= x"BF";
            when x"FF9" => q <= x"BF";
            when x"FFA" => q <= x"00";
            when x"FFB" => q <= x"00";
            when x"FFC" => q <= x"00";
            when x"FFD" => q <= x"00";
            when x"FFE" => q <= x"00";
            when x"FFF" => q <= x"00";
            when others => q <= (others => '0');
        end case;
    end process;
end RTL;
